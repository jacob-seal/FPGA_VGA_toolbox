----------------------------------------------------------------------------------
--Developed By : Jacob Seal
--sealenator@gmail.com
--07-28-2021
--filename: bitmaps_pkg.vhd
--package bitmaps_pkg
--
--********************************************************************************
--general notes:
--This package contains bitmaps that can be used to output graphics on the VGA
--      output.  
--********************************************************************************
----------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package bitmaps_pkg is

  -----------------------------------------------------------------------------
  -- Constants and bit patterns
  -----------------------------------------------------------------------------
   --array to test output of bit pattern. should output "test!" on the VGA
  type t_text_bitmap is array (0 to 14) of std_logic_vector(0 to 49);
	constant bitmap : t_text_bitmap := 
    (
        ("00000000000000000000000000000000000000000000000000"),
        ("00000000000000000000000000000000000000000000000000"),
        ("00000000000000000000000000000000000000000000000000"),
        ("00000000000000000000000000000000000000000000000000"),
        ("00000100000000000000000000000000001000000000110000"),
        ("00000100000000000000000000000000001000000000110000"),
        ("00001111000001111000000111100000011110000000110000"),
        ("00000100000011001100001000010000001000000000110000"),
        ("00000100000011111100001000000000001000000000110000"),
        ("00000100000010000000001111110000001000000000110000"),
        ("00000100000010000000000000010000001000000000000000"),
        ("00000100000010000000000000010000001000000000110000"),
        ("00000111000011111100001111100000001110000000110000"),
        ("00000000000000000000000000000000000000000000000000"),
        ("00000000000000000000000000000000000000000000000000")
    );

--     --splash page for "shitty craps" game - small version in case the large one is too many resources.
--     type t_dual_dice_bitmap is array (0 to 77) of std_logic_vector(0 to 99);
-- 	constant dual_dice_bitmap : t_dual_dice_bitmap := 
--     (
-- ("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
-- ("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
-- ("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
-- ("0000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000"),
-- ("0000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000"),
-- ("0000000000000000000000001110000000000011111111110000000000000000000000000000000000000000000000000000"),
-- ("0000000000000000000000111100001111000000000011111111110000000000000000000000000000000000000000000000"),
-- ("0000000000000000000011110000011111110000000000000011111111000000000000000000000000000000000000000000"),
-- ("0000000000000000000111000000011111110000111111000000000111000000000000000000000000000000000000000000"),
-- ("0000000000000000011100000000000111000001111111000000011111000000000000000000000000000000000000000000"),
-- ("0000000000000001110000011100000000000000111110000001110011000000000000000000000000000000000000000000"),
-- ("0000000000000111100001111111000000000000000000000011100001000000000000000000000000000000000000000000"),
-- ("0000000000001110000001111111000011111000000000001110010001000000000000000000000000000000000000000000"),
-- ("0000000000111000000000111110000111111100000000111000111001000000110000000000000000000000000000000000"),
-- ("0000000000111110000000000000000011111100000011100001111101000111111111111100000000000000000000000000"),
-- ("0000000001101111111110000000000000000000001111000001111101011110000000111111111110000000000000000000"),
-- ("0000000001100000001111111110000000000000011100000001111101111000110000000000011111111110000000000000"),
-- ("0000000001100000000000001111111111100001110000000001111111100011111110000000000000011111111100000000"),
-- ("0000000001100000000000000000000111111111000000000000111110000011111110000000000000000000011110000000"),
-- ("0000000001100000000000000000000000000110001110000000111000000001111100000000000000000000111110000000"),
-- ("0000000001100000000000000000000000000110011110000011110000000000000000000000000000000001110110000000"),
-- ("0000000001100000011000000000000000000110011111000111000000000000000000000000000000000111000110000000"),
-- ("0000000001100000111100000000000000000110011111011100000000000000000000000000000000011100000110000000"),
-- ("0000000001100001111110000000000000000010011111111000000000000000000011111100000001110000000110000000"),
-- ("0000000001100001111110000000000000000010011111100000000000000000000011111110000111000000000110000000"),
-- ("0000000001100001111110000000000000000010001111111111100000000000000011111100001110000000000110000000"),
-- ("0000000001100001111110000000000000000010000011000011111111100000000000000000111000000000000110000000"),
-- ("0000000001100000111100000000000000000010000011000000000011111111110000000011100000000000000110000000"),
-- ("0000000001100000000000000000000000000010000011000000000000000011111111111110000000000000000110000000"),
-- ("0000000001100000000000000000000000000010000011000001110000000000000000111100000000000000000110000000"),
-- ("0000000001100000000000000000000000000010000010000011111000000000000000001000000000000000000110000000"),
-- ("0000000001100000000000000000000000000010000010000011111100000011100000001100000000000000000110000000"),
-- ("0000000001100000000000000000000000000010000010000011111100000111110000001100000000000000000110000000"),
-- ("0000000001100000000000000000000000000010011110000011111100000111111000001100000000000000000110000000"),
-- ("0000000001100000000000000011100000000010111110000001111000000111111000001100000000111100000110000000"),
-- ("0000000001100000000000000111110000000010111110000000000000000111111000001100000000111100000110000000"),
-- ("0000000001100000000000001111110000000010111110000000000000000011110000001100000001111110000110000000"),
-- ("0000000001100000000000001111111000000010111110000001110000000000000000001100000001111110000110000000"),
-- ("0000000001100000000000001111111000000010011110000011111000000000000000001100000000111100000110000000"),
-- ("0000000001100000000000000111110000000010001010000011111100000011110000001100000000111100000110000000"),
-- ("0000000001100000000000000011100000000010000010000011111100000111111000001100000000000000000110000000"),
-- ("0000000001100000000000000000000000000010000010000011111100000111111000001100000000000000000110000000"),
-- ("0000000000111111000000000000000000000110000010000001111000000111111000001100000000000000000110000000"),
-- ("0000000000001111111111000000000000000110001111000000000000000111111000001100000000000000000110000000"),
-- ("0000000000000000001111111111100000000110111111000000000000000011110000001100000000000000000110000000"),
-- ("0000000000000000000000000111111111110111110011000000000000000000000000001100000000000000000110000000"),
-- ("0000000000000000000000000000000011111111000011000011111000000000000000001100000000000000001100000000"),
-- ("0000000000000000000000000000000000000000000011000011111100000011110000001100000000000000011100000000"),
-- ("0000000000000000000000000000000000000000000011000011111100000111111000001100000000000001110000000000"),
-- ("0000000000000000000000000000000000000000000011000011111100000111111000001100000000000011100000000000"),
-- ("0000000000000000000000000000000000000000000011000001111000000111111000001100000000001110000000000000"),
-- ("0000000000000000000000000000000000000000000011000000110000000011111000001100000000111000000000000000"),
-- ("0000000000000000000000000000000000000000000011111000000000000001100000001100000011110000000000000000"),
-- ("0000000000000000000000000000000000000000000000111111110000000000000000001100001111000000000000000000"),
-- ("0000000000000000000000000000000000000000000000000011111111100000000000001100111100000000000000000000"),
-- ("0000000000000000000000000000000000000000000000000000000011111111111000001111110000000000000000000000"),
-- ("0000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000"),
-- ("0000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000"),
-- ("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
-- ("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
-- ("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
-- ("0000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000"),
-- ("0000000000000001000100011000000000000000000000011100000000000000011110000011000000111100000000000000"),
-- ("0000000000010011101100011011111111111111111100011000000000111000011111000011100001110110000110000000"),
-- ("0000000011111011001111111111111101111110011100110000000111111100011011000011100000110011111110000000"),
-- ("0000000111111011001101011000011100000110011110110000000111111100011011000111110001110011111110000000"),
-- ("0000000110001011001100011000001100000110001111110000000110000000011011000111110001100011100010000000"),
-- ("0000000110000011101100011000001100000110000111110000001110000000111111000110110001100110110000000000"),
-- ("0000000011100011111000010000001000000110000111100000001110000000111111000110110001111100011000000000"),
-- ("0000000000110011001100010000001000000110000011100000001110000000111110001111111101100000001100000000"),
-- ("0000000000010011001100010000001000000110000011000000001110000110111110001111111001100000000110000000"),
-- ("0000000000011011001100010000001000000110000011000000000111001110110111001110011001000000000010000000"),
-- ("0000000000010011001100111110001000000110000011000000000011111110110011101110001101000000000110000000"),
-- ("0000000011110011001101111100001000000110000011000000000001111100110001101110001111000000111100000000"),
-- ("0000000000000011001101111000001000000100000011000000000000000000110000111100000111000000000000000000"),
-- ("0000000000000001000000000000000000000000000000000000000000000000000000011100000000000000000000000000"),
-- ("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
-- ("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000")

--     );

--splash page for "shitty craps" game
    type t_dual_dice_bitmap is array (0 to 233) of std_logic_vector(0 to 299);
	constant dual_dice_bitmap : t_dual_dice_bitmap := 
    (
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000001111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000001111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000001111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000000000000000000000000000001111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000111111100000000000000000000000000000000000000011111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000111111100000000000000001111111111111110000000000000000000000000000000000000000011111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000011111110000000000000000011111111111111111000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000111111100000000000000000111111111111111111100000000000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000011111110000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000001111111000000000000000000000111111111111111111100000000000000001111111111111000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000111111100000000000000000000000111111111111111111100000000000000111111111111111110000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000011111110000000000000000000000000011111111111111111000000000000001111111111111111111000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000011111111111000000000000000011111111111111111111000000000000000000000000011111101111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000001111110001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000111111000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000001111110000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000001111111111111000000000000000000000111111000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000111111100000000000000000111111110000000000000000000000000000000000000000000000000011100000000000000000000000011111100000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000011111110000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000111110000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000001111111000000000000000011111111111111111100000000000000000000000000000000000000000000000000000000000000000000111111100000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000011111100000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000001111110000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000001111111000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000111111100000000000000000000111111111111111111110000000000000000111111111110000000000000000000000000000000000011111100000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000011111110000000000000000000000011111111111111111100000000000000111111111111111100000000000000000000000000000000111111000000001111100000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000111111000000000000000000000000001111111111111111000000000000001111111111111111111000000000000000000000000000111111100000000111111110000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000011111110000000000000000000000000000001111111111000000000000000001111111111111111111000000000000000000000000001111110000000001111111111000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000111111100000000001111111111100000111000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000011111100000000000011111111111100000111000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000001111110000000000000011111111111110000111000000000000111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000000000011111111111111100000000000000000000111111100000000000000011111111111110000111000000000011111111000011111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000001111001111111111111111110000000000000000000000000000000000000000000000011111111100000000000000000000001111110000000000000000011111111111110000111000000001111111100000000000000011111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000001110000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000011111111111110000111000000111111110000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000001110000000000000001111111111111111100000000000000000000000000000000000000000000000000000000000000011111100000000000000000000011111111111110000111000011111110000000000000000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000001110000000000000000000001111111111111111110000000000000000000000000000000000000000000000000000001111110000000000000000000000011111111111110000111001111111000000000000000000000000000000000000000000000001111111111111111111110000000000000000000000000000000000000000000000000"),
("000000000000000000000000000001110000000000000000000000000111111111111111111111000000000000000000000000000000000000000000000111111100000000000000000000000011111111111110000111111111110000000000000000000000000000000000000000000000000000011111111111111111111110000000000000000000000000000000000000000000"),
("000000000000000000000000000001110000000000000000000000000000000011111111111111111111100000000000000000000000000000000000011111110000000000000000000000000011111111111110000111111111000000000001111111111100000000000000000000000000000000000000001111111111111111111110000000000000000000000000000000000000"),
("000000000000000000000000000001110000000000000000000000000000000000000011111111111111111111000000000000000000000000000001111111000000000000000000000000000011111111111110000111111100000000000111111111111111000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000"),
("000000000000000000000000000001110000000000000000000000000000000000000000000000111111111111111111110000000000000000000111111100000000000000000000000000000011111111111100011111100000000000011111111111111111100000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000"),
("000000000000000000000000000001110000000000000000000000000000000000000000000000000000011111111111111111111110000000011111110000000000000000000000000000000001111111111101111111000000000000011111111111111111110000000000000000000000000000000000000000000000000000000111111111111111000000000000000000000000"),
("000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000111111111111111111111111111111000000000000000000000000000000000001111111111111111100000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000000"),
("000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000111111111111110000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000"),
("000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000011111111111000000000000000000011111111111111111100000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000"),
("000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000011111000000000000000000000000000011111100000000000000000000000111111111111111000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000"),
("000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000111111100000000000000000000000001111110000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000001111111001110000000000000000000000"),
("000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000001111111110000000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100001110000000000000000000000"),
("000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000011111111111000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000001110000000000000000000000"),
("000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000011111111111100000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000001110000000000000000000000"),
("000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000111111111111100000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000001110000000000000000000000"),
("000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000111111111111100000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000001110000000000000000000000"),
("000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000111111111111100000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000001110000000000000000000000"),
("000000000000000000000000000011100000000000000000000111111000000000000000000000000000000000000000000000000000000001110000000111111111111100000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000001110000000000000000000000"),
("000000000000000000000000000011100000000000000000011111111110000000000000000000000000000000000000000000000000000001110000000111111111111100000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000001110000000000000000000000"),
("000000000000000000000000000011100000000000000000111111111111000000000000000000000000000000000000000000000000000001110000000111111111111100000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000001110000000000000000000000"),
("000000000000000000000000000011100000000000000001111111111111100000000000000000000000000000000000000000000000000001110000000111111111111100000111111100000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000111111000000000000000000001110000000000000000000000"),
("000000000000000000000000000011100000000000000011111111111111110000000000000000000000000000000000000000000000000001110000000111111111111100011111110000000000000000000000000000000000000000000000000000000000001111111111111100000000000000000000000000011111100000000000000000000001110000000000000000000000"),
("000000000000000000000000000011100000000000000011111111111111110000000000000000000000000000000000000000000000000001110000000111111111111100111111000000000000000000000000000000000000000000000000000000000000011111111111111111000000000000000000000001111110000000000000000000000001111000000000000000000000"),
("000000000000000000000000000011100000000000000111111111111111111000000000000000000000000000000000000000000000000001110000000011111111111111111100000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000111111100000000000000000000000001111000000000000000000000"),
("000000000000000000000000000111100000000000000111111111111111111000000000000000000000000000000000000000000000000001110000000011111111111111111000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000011111100000000000000000000000000001111000000000000000000000"),
("000000000000000000000000000111100000000000000111111111111111111000000000000000000000000000000000000000000000000001110000000001111111111111100000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000111111000000000000000000000000000001111000000000000000000000"),
("000000000000000000000000000111100000000000000111111111111111111000000000000000000000000000000000000000000000000001110000000001111111111111111111000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000011111100000000000000000000000000000001111000000000000000000000"),
("000000000000000000000000000111100000000000000111111111111111111000000000000000000000000000000000000000000000000001110000000000111111111111111111111100000000000000000000000000000000000000000000000000000000011111111111111111000000000000001111110000000000000000000000000000000001111000000000000000000000"),
("000000000000000000000000000111100000000000000111111111111111111000000000000000000000000000000000000000000000000001110000000000000000011100111111111111111100000000000000000000000000000000000000000000000000000111111111111000000000000000111111100000000000000000000000000000000001111000000000000000000000"),
("000000000000000000000000000111100000000000000011111111111111110000000000000000000000000000000000000000000000000001110000000000000000011100000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000001111000000000000000000000"),
("000000000000000000000000000111100000000000000011111111111111110000000000000000000000000000000000000000000000000001110000000000000000011100000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000001111000000000000000000000"),
("000000000000000000000000000111100000000000000001111111111111100000000000000000000000000000000000000000000000000001110000000000000000111100000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000001111000000000000000000000"),
("000000000000000000000000000111100000000000000000111111111111100000000000000000000000000000000000000000000000000001110000000000000000111100000000000000000000000011111111111111111100000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000001111000000000000000000000"),
("000000000000000000000000000111100000000000000000011111111110000000000000000000000000000000000000000000000000000001110000000000000000111100000000000000000000000000000001111111111111111110000000000000000000000000000000000000000111111000000000000000000000000000000000000000000001111000000000000000000000"),
("000000000000000000000000000111100000000000000000001111111100000000000000000000000000000000000000000000000000000001110000000000000000111100000000000000000000000000000000000001111111111111111111100000000000000000000000000000011111110000000000000000000000000000000000000000000001111000000000000000000000"),
("000000000000000000000000000111100000000000000000000001110000000000000000000000000000000000000000000000000000000001110000000000000000111100000000000000000000000000000000000000000011111111111111111111111000000000000000000001111111000000000000000000000000000000000000000000000001111000000000000000000000"),
("000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000111100000000000000000000000000000000000000000000000001111111111111111111110000000000000011111100000000000000000000000000000000000000000000000001111000000000000000000000"),
("000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000111100000000000000000000000000000000000000000000000000000000011111111111111111111110001111110000000000000000000000000000000000000000000000000001111000000000000000000000"),
("000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000111100000000000000000000000000000000000000000000000000000000000000000111111111111111111111000000000000000000000000000000000000000000000000000001111000000000000000000000"),
("000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000001111000000000000000000000"),
("000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000111100000000000000000000111000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000001111000000000000000000000"),
("000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000111100000000000000000011111111000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000001111000000000000000000000"),
("000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000111100000000000000001111111111110000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000001111000000000000000000000"),
("000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000111100000000000000011111111111111000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000001111000000000000000000000"),
("000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000111100000000000000011111111111111000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000001111000000000000000000000"),
("000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000111000000000000000111111111111111100000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000001111000000000000000000000"),
("000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000111000000000000000111111111111111110000000000000000000000010000000000000000000000000011100000000000000000000000000000000000000000000000000000001111000000000000000000000"),
("000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000111000000000000000111111111111111110000000000000000000011111111100000000000000000000011100000000000000000000000000000000000000000000000000000001111000000000000000000000"),
("000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000111000000000000000111111111111111110000000000000000001111111111110000000000000000000011100000000000000000000000000000000000000000000000000000001111000000000000000000000"),
("000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000111000000000000000111111111111111110000000000000000011111111111111000000000000000000011100000000000000000000000000000000000000000000000000000001111000000000000000000000"),
("000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000011100111000000000000000111111111111111110000000000000000011111111111111100000000000000000011100000000000000000000000000000000000000000000000000000001111000000000000000000000"),
("000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000001111110111000000000000000111111111111111110000000000000000011111111111111100000000000000000011100000000000000000000000000000000000000000000000000000001111000000000000000000000"),
("000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000011111111111000000000000000011111111111111110000000000000000111111111111111110000000000000000011100000000000000000000000000000000000000000000000000000001111000000000000000000000"),
("000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000111111111111000000000000000011111111111111100000000000000000111111111111111110000000000000000011100000000000000000000000000000011110000000000000000000001111000000000000000000000"),
("000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000111111111111000000000000000001111111111111000000000000000000111111111111111111000000000000000011100000000000000000000000000001111111100000000000000000001111000000000000000000000"),
("000000000000000000000000000011100000000000000000000000000000000000000000000000000111000000000000000000000000000001110000001111111111111000000000000000000111111111110000000000000000000111111111111111111000000000000000011100000000000000000000000000011111111110000000000000000001111000000000000000000000"),
("000000000000000000000000000011100000000000000000000000000000000000000000000000111111110000000000000000000000000001110000001111111111111000000000000000000001111111100000000000000000000011111111111111111000000000000000011100000000000000000000000000011111111110000000000000000001111000000000000000000000"),
("000000000000000000000000000011100000000000000000000000000000000000000000000001111111111100000000000000000000000001110000001111111111111000000000000000000000000000000000000000000000000011111111111111110000000000000000011100000000000000000000000000111111111111000000000000000001111000000000000000000000"),
("000000000000000000000000000011110000000000000000000000000000000000000000000011111111111110000000000000000000000001110000011111111111111000000000000000000000000000000000000000000000000011111111111111110000000000000000011100000000000000000000000000111111111111100000000000000001111000000000000000000000"),
("000000000000000000000000000011110000000000000000000000000000000000000000000111111111111111000000000000000000000001110000011111111111111000000000000000000000000000000000000000000000000001111111111111100000000000000000011100000000000000000000000001111111111111100000000000000001111000000000000000000000"),
("000000000000000000000000000011110000000000000000000000000000000000000000001111111111111111000000000000000000000001110000011111111111111000000000000000000000000000000000000000000000000000111111111111100000000000000000011100000000000000000000000001111111111111100000000000000001111000000000000000000000"),
("000000000000000000000000000011110000000000000000000000000000000000000000001111111111111111100000000000000000000001110000011111111111111000000000000000000000000000000000000000000000000000011111111111000000000000000000011100000000000000000000000001111111111111100000000000000001110000000000000000000000"),
("000000000000000000000000000011110000000000000000000000000000000000000000001111111111111111100000000000000000000001110000001111111111111000000000000000000000000000000000000000000000000000000011111000000000000000000000011100000000000000000000000001111111111111100000000000000001110000000000000000000000"),
("000000000000000000000000000001110000000000000000000000000000000000000000011111111111111111100000000000000000000001110000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000001111111111111100000000000000001110000000000000000000000"),
("000000000000000000000000000001110000000000000000000000000000000000000000011111111111111111100000000000000000000001110000001111111111111000000000000000000011111111000000000000000000000000000000000000000000000000000000001100000000000000000000000001111111111111100000000000000001110000000000000000000000"),
("000000000000000000000000000001110000000000000000000000000000000000000000011111111111111111100000000000000000000001110000001111111111111000000000000000001111111111100000000000000000000000000000000000000000000000000000001110000000000000000000000001111111111111100000000000000001110000000000000000000000"),
("000000000000000000000000000001110000000000000000000000000000000000000000001111111111111111100000000000000000000001110000000111111111111000000000000000011111111111110000000000000000000000000000000000000000000000000000001110000000000000000000000000111111111111100000000000000001110000000000000000000000"),
("000000000000000000000000000001110000000000000000000000000000000000000000001111111111111111100000000000000000000001110000000111111111111000000000000000011111111111111000000000000000000000000000000000000000000000000000001110000000000000000000000000111111111111000000000000000001110000000000000000000000"),
("000000000000000000000000000001110000000000000000000000000000000000000000001111111111111111100000000000000000000001110000000011111111111000000000000000111111111111111100000000000000000000000000000000000000000000000000001110000000000000000000000000111111111111000000000000000001110000000000000000000000"),
("000000000000000000000000000001110000000000000000000000000000000000000000000111111111111111000000000000000000000001110000000001111110111000000000000000111111111111111110000000000000000000000111100000000000000000000000001110000000000000000000000000011111111110000000000000000001110000000000000000000000"),
("000000000000000000000000000001110000000000000000000000000000000000000000000111111111111110000000000000000000000001110000000000000000111000000000000000111111111111111110000000000000000000011111111000000000000000000000001110000000000000000000000000011111111110000000000000000001110000000000000000000000"),
("000000000000000000000000000001110000000000000000000000000000000000000000000011111111111100000000000000000000000001110000000000000000111000000000000000111111111111111110000000000000000000111111111110000000000000000000001110000000000000000000000000001111111100000000000000000001110000000000000000000000"),
("000000000000000000000000000001110000000000000000000000000000000000000000000001111111111000000000000000000000000001110000000000000000111000000000000000111111111111111110000000000000000001111111111111000000000000000000001110000000000000000000000000000001110000000000000000000001110000000000000000000000"),
("000000000000000000000000000001110000000000000000000000000000000000000000000000011111110000000000000000000000000001110000000000000000111000000000000000111111111111111110000000000000000011111111111111100000000000000000001110000000000000000000000000000000000000000000000000000001110000000000000000000000"),
("000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000111000000000000000111111111111111110000000000000000011111111111111100000000000000000001110000000000000000000000000000000000000000000000000000001110000000000000000000000"),
("000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000111000000000000000011111111111111110000000000000000111111111111111110000000000000000001110000000000000000000000000000000000000000000000000000001110000000000000000000000"),
("000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000111000000000000000011111111111111100000000000000000111111111111111110000000000000000001110000000000000000000000000000000000000000000000000000001110000000000000000000000"),
("000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000111000000000000000001111111111111000000000000000000111111111111111111000000000000000001110000000000000000000000000000000000000000000000000000001110000000000000000000000"),
("000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000111000000000000000000111111111110000000000000000000111111111111111111000000000000000001110000000000000000000000000000000000000000000000000000001110000000000000000000000"),
("000000000000000000000000000000111111111110000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000111100000000000000000001111111100000000000000000000011111111111111111000000000000000001110000000000000000000000000000000000000000000000000000001110000000000000000000000"),
("000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000001110000000000000000111100000000000000000000000000000000000000000000000011111111111111110000000000000000001110000000000000000000000000000000000000000000000000000001110000000000000000000000"),
("000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000000000000001110000000000000011111100000000000000000000000000000000000000000000000011111111111111110000000000000000001110000000000000000000000000000000000000000000000000000001110000000000000000000000"),
("000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000000000001110000000000000111111100000000000000000000000000000000000000000000000001111111111111100000000000000000001110000000000000000000000000000000000000000000000000000011110000000000000000000000"),
("000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000001110000000000011111111100000000000000000000000000000000000000000000000000111111111111100000000000000000001110000000000000000000000000000000000000000000000000000011110000000000000000000000"),
("000000000000000000000000000000000000000000000000000011111111111111111111100000000000000000000000000000000000000001110000000001111111111100000000000000000000000000000000000000000000000000011111111111000000000000000000001110000000000000000000000000000000000000000000000000000011110000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000111111111111111111111000000000000000000000000000000001110000000111111100111100000000000000000000000000000000000000000000000000000111111100000000000000000000001110000000000000000000000000000000000000000000000000000011110000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000011111111111111111111110000000000000000000000001110000011111110000111100000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000011110000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111000000000000000001110011111111100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000011110000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111110000000001111111111100000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000011100000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111100001111111110000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000011100000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111000000000000111100000000000000000011111111000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000111100000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111000000000000000111100000000000000001111111111110000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000001111000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000011100000000000000011111111111111000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000011111000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000011111111111111100000000000000000000001111111000000000000000000000001110000000000000000000000000000000000000000000000001111110000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000111111111111111100000000000000000000111111111110000000000000000000001110000000000000000000000000000000000000000000000011111100000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000111111111111111110000000000000000001111111111111000000000000000000001110000000000000000000000000000000000000000000001111110000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000111111111111111110000000000000000011111111111111100000000000000000001110000000000000000000000000000000000000000000011111100000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000111111111111111110000000000000000011111111111111100000000000000000001110000000000000000000000000000000000000000001111110000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000111111111111111110000000000000000011111111111111110000000000000000001110000000000000000000000000000000000000000111111100000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000111111111111111110000000000000000111111111111111110000000000000000001110000000000000000000000000000000000000001111110000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000111111111111111110000000000000000111111111111111111000000000000000001110000000000000000000000000000000000000111111100000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000011111111111111110000000000000000111111111111111111000000000000000001110000000000000000000000000000000000011111110000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000001111111111111100000000000000000111111111111111111000000000000000001110000000000000000000000000000000001111111100000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000111111111111000000000000000000011111111111111110000000000000000001100000000000000000000000000000000011111100000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000011111111110000000000000000000011111111111111110000000000000000011100000000000000000000000000000001111111000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000111111000000000000000000000001111111111111100000000000000000011100000000000000000000000000000111111100000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000111111111111100000000000000000011100000000000000000000000000011111111000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000011111111111000000000000000000011100000000000000000000000000111111100000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000001111111110000000000000000000011100000000000000000000000011111110000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000100000000000000000000000011100000000000000000000001111111000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000111111100000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000011100000000000000000011111110000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000000000000000000011100000000000000001111111000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000011100000000000000111111110000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000000011100000000000011111110000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000011100000000001111111000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111000000000000000000000000000000000000011100000001111111110000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000000011100000011111111000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111000000000000000000000000011100001111111000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111100000000000000011100111111100000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000010000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000110000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000001110000000000111110000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000111111110000000000000000011110000000000000000000111111111111000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000011111100000001110000000000111110000000000000000000000111100000000000000000011110011111000000000000011111000000000000000000000000000000000000000000000000011111111111100000000000000111111000000000000000001111111111111100000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000011111100000001110000000000111110000000111111111111111111111111111111111111111111111111110000000000111110000000000000000000000000000000000000000000000000111111111111110000000000000111111100000000000000001111110001111110000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000011111110000001110000000000111110000011111111111111111111111111111111111111111111111111110000000000111100000000000000000000000000000011111100000000000000111111111111110000000000000011111100000000000000001111110000011111000000000000000000000000000000000000000"),
("000000000000000000000000000000011111000000011111100000011110000000000111110000011111111111111111111111111111111111111111111111111111000000001111100000000000000000000000000011111111111000000000000111111001111111000000000000011111100000000000000001111110000001111000000000000111110000000000000000000000"),
("000000000000000000000000001111111111100000011111100000011100011110000111111111111111111111111000000011111111111111100000001111111111000000001111000000000000000000000000011111111111111000000000000111110000111111000000000000111111110000000000000001111110000001111000000011111111110000000000000000000000"),
("000000000000000000000000011111111111100000011111100000011100111111111111111111111111111111111100000001111111111111100000000111111111000000011111000000000000000000000001111111111111111100000000000111110000111111000000000000111111111000000000000001111110000000111100001111111111111000000000000000000000"),
("000000000000000000000000111111111111110000011111000000011100111111111111110000000111111111111100000000111111111111110000000011111111000000011110000000000000000000000011111111111111111110000000000111110000111111100000000001111111111000000000000001111100000000111100011111111111111000000000000000000000"),
("000000000000000000000001111111111111110000011111000000011100011111000111100000000000000001111110000000000000000111110000000001111111100000111110000000000000000000000111111111111111111110000000000111110001111111100000000001111111111100000000000001111100000000111100111111111111111000000000000000000000"),
("000000000000000000000011111100000111110000011111000000011100000000000111100000000000000001111110000000000000000111110000000001111111100000111110000000000000000000000111111111000011111100000000000111110000111111100000000001111111111100000000000111111100000000111101111111000011111100000000000000000000"),
("000000000000000000000111111000000011110000011110000000011100000000000111100000000000000001111100000000000000000111110000000000111111100000111110000000000000000000000111111100000000010000000000000111100001111111100000000001111111111100000000000011111100000000111101111100000001111100000000000000000000"),
("000000000000000000000111110000000001110000011110000000011100000000000111100000000000000001111100000000000000000111110000000000011111110000111110000000000000000000000111111000000000000000000000000111100001111111100000000001111001111110000000000001111100000000111101111100000000111100000000000000000000"),
("000000000000000000000111110000000000000000011110000000111100000000000111100000000000000000111100000000000000000011110000000000001111110001111110000000000000000000001111111000000000000000000000001111100001111111100000000001111001111110000000000011111100000000111101111000000000000000000000000000000000"),
("000000000000000000000111110000000000000000011110000000111100000000000111100000000000000000111100000000000000000011110000000000000111111001111110000000000000000000001111110000000000000000000000001111100001111111000000000011111001111110000000000011111000000000111101111000000000000000000000000000000000"),
("000000000000000000000011110000000000000000011110000000111100000000000111100000000000000000111100000000000000000011110000000000000011111011111100000000000000000000001111110000000000000000000000001111000001111111000000000011111001111110000000000011111000000001111001111100000000000000000000000000000000"),
("000000000000000000000011111000000000000000111111000000111100000000000111100000000000000000111100000000000000000011110000000000000111111111111100000000000000000000011111110000000000000000000000001111001111111111000000000011111000111111000000000011111000000001111001111110000000000000000000000000000000"),
("000000000000000000000001111100000000000001111111111111111100000000000111100000000000000000111100000000000000000111110000000000000111111111111000000000000000000000011111100000000000000000000000001111111111111111000000000011111000111111000000000011111011100011110000111111000000000000000000000000000000"),
("000000000000000000000000111111000000000001111111111111111100000000000111100000000000000000111100000000000000000111100000000000000111111111110000000000000000000000011111100000000000000000000000001111111111111110000000000011111000111111000000000011111011111111100000011111100000000000000000000000000000"),
("000000000000000000000000001111100000000001111111111111111100000000000111100000000000000000111100000000000000000111100000000000000011111111110000000000000000000000011111100000000000000000000000001111111111111000000000000011111000111111000000000011111001111110000000000111111000000000000000000000000000"),
("000000000000000000000000000111111000000000111110000011111100000000000111100000000000000000111000000000000000000011100000000000000001111111100000000000000000000000011111100000000000000000000000001111111111110000000000001111111110011111100000000011110000000000000000000001111100000000000000000000000000"),
("000000000000000000000000000001111100000000011110000000111100000000000111100000000000000000111000000000000000000011100000000000000001111111100000000000000000000000011111100000000000000000000000001111111111110000000000001111111111111111100000000011110000000000000000000000111110000000000000000000000000"),
("000000000000000000000000000000111110000000011110000000111100000000000111100000000000000000111000000000000000000011100000000000000000111111100000000000000000000000011111100000000000000000000000011111111111110000000000001111111111111111111111000011110000000000000000000000001111000000000000000000000000"),
("000000000000000000000000000000011110000000011110000000111100000000000111100000000000000000111000000000000000000111100000000000000000111111100000000000000000000000011111100000000000000000000000011110011111111000000000001111111111111111111111000011110000000000000000000000000111100000000000000000000000"),
("000000000000000000000000000000001111000000011110000001111100000000000111100000000000000000111000000000000000000111100000000000000000111111000000000000000000000000001111100000000000000000111000011110001111111000000000011111111111111111111100000111110000000000000000000000000011100000000000000000000000"),
("000000000000000000000000000000000111000000011110000000111100000000000111100000000000000000111000000000000000000011100000000000000000111111000000000000000000000000001111110000000000000011111000011110001111111100000000011111111111111111110000000111100000000000000000000000000011110000000000000000000000"),
("000000000000000000000000000000000111100000011110000001111100000000000111100000000000000000111000000000000000000011100000000000000000111111000000000000000000000000001111110000000000000111111000011110100111111100000000011111111110000111110000000111100000000000000000000000000001110000000000000000000000"),
("000000000000000000000000000000000011100000011110000001111100000000000111100000000000000000111000000000000000000011100000000000000000111111000000000000000000000000000111111000000000001111111000011110000011111110000000011111111100000011111000000111100000000000000000000000000001110000000000000000000000"),
("000000000000000000000000000000000011100000011110000000111100000000000111100000000000000000111000000000000000000011100000000000000000011111000000000000000000000000000011111100000000001111110000011100000001111110000000001111111000000001111000000111100000000000000000000000000001111000000000000000000000"),
("000000000000000000000000000000000011100000011100000000111100000000000111100000000000000000111000000000000000000011100000000000000000011110000000000000000000000000000011111110000000011111110000011100000000111111000000001111100000000001111000000111000000000000000000000000000000111000000000000000000000"),
("000000000000000000000000000000000011100000011100000000111100000000000111111100011100000000111000000000000000000011100000000000000000011110000000000000000000000000000001111111000001111111110000111100000000111111000000001111100000000000111100001111000000000000000000000000000001110000000000000000000000"),
("000000000000000000000000000000000111100000011100000000111100000000111111111111101000000000111000000000000000000011100000000000000000111110000000000000000000000000000000011111111111111111100000111100000000011111100000001111100000000000011100001111000000000000000000000000000001110000000000000000000000"),
("000000000000000000000000000000000111000000011100000000111100000011111111111111111000000000111000000000000000000011100000000000000000111110000000000000000000000000000000001111111111111111000000111100000000001111100000011111100000000000011110001110000000000000000000000000000001110000000000000000000000"),
("000000000000000000000000000000000111000000011100000000111110000011111111111111110000000000111000000000000000000011100000000000000000111100000000000000000000000000000000000111111111111110000000111100000000000111110001111111100000000000011110001110000000000000000000000000000011100000000000000000000000"),
("000000000000000000000000111000011110000000011100000000111110000111111111111000000000000000111000000000000000000011100000000000000000111100000000000000000000000000000000000001111111111100000000111100000000000011110000111111100000000000001110001110000000000000000000001100000111000000000000000000000000"),
("000000000000000000000000111111111100000000011100000000111110000111111111100000000000000000011000000000000000000011100000000000000000111100000000000000000000000000000000000000011111111000000000111100000000000001111001111111100000000000001111001110000000000000000000001111111110000000000000000000000000"),
("000000000000000000000000001111100000000000011100000000011111000111111111100000000000000000011000000000000000000011100000000000000000011100000000000000000000000000000000000000000000000000000000111100000000000001111001111111100000000000000111001110000000000000000000000011110000000000000000000000000000"),
("000000000000000000000000000000000000000000011100000000001111000011111111100000000000000000011000000000000000000011100000000000000000011100000000000000000000000000000000000000000000000000000000011110000000000000111101111111000000000000000111101110000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000011100000000000110000001111100000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000011100000000000000011111111111000000000000000011101110000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000")



    );


    --define array to hold large dice bitmaps
    type t_large_dice_bitmap is array (0 to 149) of std_logic_vector(0 to 146);
	
    --dice number 1
    constant large_dice_bitmap_1 : t_large_dice_bitmap := 
    (
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000011111111111000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000001111111111111110000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000011111111111111111000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000001111111111111111111110000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000011111111111111111111110000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000001111111111111111111110000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000011111111111111111000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000001111111111111110000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000111111111111100000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000111111100000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000"),
("000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000")

);

     --dice number 2
	constant large_dice_bitmap_2 : t_large_dice_bitmap := 
    (
        ("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000011111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000001111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000001111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000001111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000001111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000001111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000001111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111100000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111110000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111110000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111110000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111100000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000"),
("000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000")

    );

     --dice number 3
	constant large_dice_bitmap_3 : t_large_dice_bitmap := 
    (
        ("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000001111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000011111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000011111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000001111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000001111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000011111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000011111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000001111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000011111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000111111111111100000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000011111111111111111111110000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000001111111111111111111111111110000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000001111111111111111111111111110000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000011111111111111111111110000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000001111111111111111111110000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000111111111111100000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111100000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111100000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111100000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111100000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111110000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111100000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111100000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111110000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000"),
("000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000")

    );

     --dice number 4
	constant large_dice_bitmap_4 : t_large_dice_bitmap := 
    (
        ("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000111111100000000000000000000000000000000000000000000000000000000011111110000000000000000000000000001000000000"),
("000000000001000000000000000000000000011111111111100000000000000000000000000000000000000000000000000011111111111100000000000000000000000001000000000"),
("000000000001000000000000000000000001111111111111111000000000000000000000000000000000000000000000001111111111111111000000000000000000000001000000000"),
("000000000001000000000000000000000011111111111111111100000000000000000000000000000000000000000000011111111111111111100000000000000000000001000000000"),
("000000000001000000000000000000000111111111111111111110000000000000000000000000000000000000000000111111111111111111110000000000000000000001000000000"),
("000000000001000000000000000000001111111111111111111111000000000000000000000000000000000000000001111111111111111111111000000000000000000001000000000"),
("000000000001000000000000000000011111111111111111111111000000000000000000000000000000000000000001111111111111111111111100000000000000000001000000000"),
("000000000001000000000000000000011111111111111111111111100000000000000000000000000000000000000011111111111111111111111100000000000000000001000000000"),
("000000000001000000000000000000111111111111111111111111100000000000000000000000000000000000000011111111111111111111111110000000000000000001000000000"),
("000000000001000000000000000000111111111111111111111111100000000000000000000000000000000000000111111111111111111111111110000000000000000001000000000"),
("000000000001000000000000000000111111111111111111111111110000000000000000000000000000000000000111111111111111111111111110000000000000000001000000000"),
("000000000001000000000000000000111111111111111111111111110000000000000000000000000000000000000111111111111111111111111110000000000000000001000000000"),
("000000000001000000000000000000111111111111111111111111110000000000000000000000000000000000000111111111111111111111111110000000000000000001000000000"),
("000000000001000000000000000000111111111111111111111111110000000000000000000000000000000000000111111111111111111111111110000000000000000001000000000"),
("000000000001000000000000000000111111111111111111111111110000000000000000000000000000000000000111111111111111111111111110000000000000000001000000000"),
("000000000001000000000000000000111111111111111111111111110000000000000000000000000000000000000111111111111111111111111110000000000000000001000000000"),
("000000000001000000000000000000111111111111111111111111100000000000000000000000000000000000000011111111111111111111111110000000000000000001000000000"),
("000000000001000000000000000000011111111111111111111111100000000000000000000000000000000000000011111111111111111111111100000000000000000001000000000"),
("000000000001000000000000000000011111111111111111111111000000000000000000000000000000000000000001111111111111111111111100000000000000000001000000000"),
("000000000001000000000000000000001111111111111111111111000000000000000000000000000000000000000001111111111111111111111000000000000000000001000000000"),
("000000000001000000000000000000000111111111111111111110000000000000000000000000000000000000000000111111111111111111110000000000000000000001000000000"),
("000000000001000000000000000000000011111111111111111100000000000000000000000000000000000000000000011111111111111111100000000000000000000001000000000"),
("000000000001000000000000000000000001111111111111111000000000000000000000000000000000000000000000001111111111111111000000000000000000000001000000000"),
("000000000001000000000000000000000000011111111111100000000000000000000000000000000000000000000000000011111111111100000000000000000000000001000000000"),
("000000000001000000000000000000000000000111111100000000000000000000000000000000000000000000000000000000011111110000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000001000000000"),
("000000000001000000000000000000000000011111111111000000000000000000000000000000000000000000000000000001111111111100000000000000000000000001000000000"),
("000000000001000000000000000000000001111111111111110000000000000000000000000000000000000000000000000111111111111110000000000000000000000001000000000"),
("000000000001000000000000000000000011111111111111111000000000000000000000000000000000000000000000001111111111111111100000000000000000000001000000000"),
("000000000001000000000000000000000111111111111111111100000000000000000000000000000000000000000000011111111111111111110000000000000000000001000000000"),
("000000000001000000000000000000001111111111111111111110000000000000000000000000000000000000000000111111111111111111111000000000000000000001000000000"),
("000000000001000000000000000000011111111111111111111111000000000000000000000000000000000000000001111111111111111111111000000000000000000001000000000"),
("000000000001000000000000000000011111111111111111111111100000000000000000000000000000000000000011111111111111111111111100000000000000000001000000000"),
("000000000001000000000000000000111111111111111111111111100000000000000000000000000000000000000011111111111111111111111110000000000000000001000000000"),
("000000000001000000000000000000111111111111111111111111100000000000000000000000000000000000000011111111111111111111111110000000000000000001000000000"),
("000000000001000000000000000000111111111111111111111111110000000000000000000000000000000000000111111111111111111111111110000000000000000001000000000"),
("000000000001000000000000000000111111111111111111111111110000000000000000000000000000000000000111111111111111111111111110000000000000000001000000000"),
("000000000001000000000000000000111111111111111111111111110000000000000000000000000000000000000111111111111111111111111110000000000000000001000000000"),
("000000000001000000000000000000111111111111111111111111110000000000000000000000000000000000000111111111111111111111111110000000000000000001000000000"),
("000000000001000000000000000000111111111111111111111111110000000000000000000000000000000000000111111111111111111111111110000000000000000001000000000"),
("000000000001000000000000000000111111111111111111111111110000000000000000000000000000000000000111111111111111111111111110000000000000000001000000000"),
("000000000001000000000000000000111111111111111111111111100000000000000000000000000000000000000011111111111111111111111110000000000000000001000000000"),
("000000000001000000000000000000011111111111111111111111100000000000000000000000000000000000000011111111111111111111111100000000000000000001000000000"),
("000000000001000000000000000000011111111111111111111111000000000000000000000000000000000000000011111111111111111111111100000000000000000001000000000"),
("000000000001000000000000000000001111111111111111111111000000000000000000000000000000000000000001111111111111111111111000000000000000000001000000000"),
("000000000001000000000000000000001111111111111111111110000000000000000000000000000000000000000000111111111111111111111000000000000000000001000000000"),
("000000000001000000000000000000000111111111111111111100000000000000000000000000000000000000000000011111111111111111110000000000000000000001000000000"),
("000000000001000000000000000000000011111111111111111000000000000000000000000000000000000000000000001111111111111111100000000000000000000001000000000"),
("000000000001000000000000000000000000111111111111110000000000000000000000000000000000000000000000000111111111111110000000000000000000000001000000000"),
("000000000001000000000000000000000000001111111111000000000000000000000000000000000000000000000000000001111111111000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000"),
("000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000")

    );

     --dice number 5
	constant large_dice_bitmap_5 : t_large_dice_bitmap := 
    (
        ("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000001111000000000000000000000000000000000000000000000000000000001111000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000001111111111000000000000000000000000000000000000000000000000001111111111000000000000000000000000010000000000000"),
("000000000000100000000000000000000000111111111111110000000000000000000000000000000000000000000000111111111111110000000000000000000000010000000000000"),
("000000000000100000000000000000000001111111111111111000000000000000000000000000000000000000000001111111111111111000000000000000000000010000000000000"),
("000000000000100000000000000000000011111111111111111100000000000000000000000000000000000000000011111111111111111100000000000000000000010000000000000"),
("000000000000100000000000000000000111111111111111111110000000000000000000000000000000000000000111111111111111111110000000000000000000010000000000000"),
("000000000000100000000000000000001111111111111111111111000000000000000000000000000000000000000111111111111111111111000000000000000000010000000000000"),
("000000000000100000000000000000001111111111111111111111000000000000000000000000000000000000001111111111111111111111000000000000000000010000000000000"),
("000000000000100000000000000000011111111111111111111111100000000000000000000000000000000000001111111111111111111111100000000000000000010000000000000"),
("000000000000100000000000000000011111111111111111111111100000000000000000000000000000000000011111111111111111111111100000000000000000010000000000000"),
("000000000000100000000000000000011111111111111111111111100000000000000000000000000000000000011111111111111111111111100000000000000000010000000000000"),
("000000000000100000000000000000011111111111111111111111100000000000000000000000000000000000011111111111111111111111110000000000000000010000000000000"),
("000000000000100000000000000000011111111111111111111111100000000000000000000000000000000000011111111111111111111111110000000000000000010000000000000"),
("000000000000100000000000000000011111111111111111111111100000000000000000000000000000000000011111111111111111111111110000000000000000010000000000000"),
("000000000000100000000000000000011111111111111111111111100000000000000000000000000000000000011111111111111111111111110000000000000000010000000000000"),
("000000000000100000000000000000011111111111111111111111100000000000000000000000000000000000011111111111111111111111110000000000000000010000000000000"),
("000000000000100000000000000000011111111111111111111111100000000000000000000000000000000000011111111111111111111111100000000000000000010000000000000"),
("000000000000100000000000000000011111111111111111111111100000000000000000000000000000000000001111111111111111111111100000000000000000010000000000000"),
("000000000000100000000000000000001111111111111111111111000000000000000000000000000000000000001111111111111111111111100000000000000000010000000000000"),
("000000000000100000000000000000001111111111111111111111000000000000000000000000000000000000001111111111111111111111000000000000000000010000000000000"),
("000000000000100000000000000000000111111111111111111110000000000000000000000000000000000000000111111111111111111110000000000000000000010000000000000"),
("000000000000100000000000000000000011111111111111111100000000000000000000000000000000000000000011111111111111111110000000000000000000010000000000000"),
("000000000000100000000000000000000001111111111111111000000000000000000000000000000000000000000001111111111111111100000000000000000000010000000000000"),
("000000000000100000000000000000000000111111111111110000000000000000000000000000000000000000000000111111111111111000000000000000000000010000000000000"),
("000000000000100000000000000000000000011111111111100000000000000000000000000000000000000000000000001111111111100000000000000000000000010000000000000"),
("000000000000100000000000000000000000000011111100000000000000000000000000000000000000000000000000000011111100000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000001111111111100000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000011111111111111111100000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000001111111111111111111111000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000001111111111111111111111000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000011111111111111111111111110000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000011111111111111111111111110000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000011111111111111111111111110000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000011111111111111111111111110000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000001111111111111111111111000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000001111111111111111111111000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000011111111111111111100000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000001111111111100000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000011111100000000000000000000000000000000000000000000000000000011111110000000000000000000000000010000000000000"),
("000000000000100000000000000000000000011111111111100000000000000000000000000000000000000000000000001111111111100000000000000000000000010000000000000"),
("000000000000100000000000000000000000111111111111110000000000000000000000000000000000000000000000111111111111111000000000000000000000010000000000000"),
("000000000000100000000000000000000001111111111111111100000000000000000000000000000000000000000001111111111111111100000000000000000000010000000000000"),
("000000000000100000000000000000000011111111111111111100000000000000000000000000000000000000000011111111111111111110000000000000000000010000000000000"),
("000000000000100000000000000000000111111111111111111110000000000000000000000000000000000000000111111111111111111110000000000000000000010000000000000"),
("000000000000100000000000000000001111111111111111111111000000000000000000000000000000000000001111111111111111111111000000000000000000010000000000000"),
("000000000000100000000000000000001111111111111111111111000000000000000000000000000000000000001111111111111111111111100000000000000000010000000000000"),
("000000000000100000000000000000011111111111111111111111100000000000000000000000000000000000001111111111111111111111100000000000000000010000000000000"),
("000000000000100000000000000000011111111111111111111111100000000000000000000000000000000000011111111111111111111111100000000000000000010000000000000"),
("000000000000100000000000000000011111111111111111111111100000000000000000000000000000000000011111111111111111111111110000000000000000010000000000000"),
("000000000000100000000000000000011111111111111111111111100000000000000000000000000000000000011111111111111111111111110000000000000000010000000000000"),
("000000000000100000000000000000011111111111111111111111100000000000000000000000000000000000011111111111111111111111110000000000000000010000000000000"),
("000000000000100000000000000000011111111111111111111111100000000000000000000000000000000000011111111111111111111111110000000000000000010000000000000"),
("000000000000100000000000000000011111111111111111111111100000000000000000000000000000000000011111111111111111111111110000000000000000010000000000000"),
("000000000000100000000000000000011111111111111111111111100000000000000000000000000000000000011111111111111111111111100000000000000000010000000000000"),
("000000000000100000000000000000011111111111111111111111100000000000000000000000000000000000011111111111111111111111100000000000000000010000000000000"),
("000000000000100000000000000000011111111111111111111111100000000000000000000000000000000000001111111111111111111111100000000000000000010000000000000"),
("000000000000100000000000000000001111111111111111111111000000000000000000000000000000000000001111111111111111111111000000000000000000010000000000000"),
("000000000000100000000000000000001111111111111111111111000000000000000000000000000000000000000111111111111111111111000000000000000000010000000000000"),
("000000000000100000000000000000000111111111111111111110000000000000000000000000000000000000000111111111111111111110000000000000000000010000000000000"),
("000000000000100000000000000000000011111111111111111100000000000000000000000000000000000000000011111111111111111100000000000000000000010000000000000"),
("000000000000100000000000000000000001111111111111111000000000000000000000000000000000000000000001111111111111111000000000000000000000010000000000000"),
("000000000000100000000000000000000000111111111111110000000000000000000000000000000000000000000000111111111111110000000000000000000000010000000000000"),
("000000000000100000000000000000000000001111111111000000000000000000000000000000000000000000000000001111111111000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000001111000000000000000000000000000000000000000000000000000000001111000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000"),
("000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000")

    );

     --dice number 6
	constant large_dice_bitmap_6 : t_large_dice_bitmap := 
    (
        ("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000011111110000000000000000000000000000000000000000000000000000011111110000000000000000000000000001000000000000"),
("000000000000100000000000000000000000011111111111100000000000000000000000000000000000000000000000001111111111110000000000000000000000001000000000000"),
("000000000000100000000000000000000000111111111111111000000000000000000000000000000000000000000000111111111111111000000000000000000000001000000000000"),
("000000000000100000000000000000000001111111111111111100000000000000000000000000000000000000000001111111111111111100000000000000000000001000000000000"),
("000000000000100000000000000000000011111111111111111110000000000000000000000000000000000000000011111111111111111110000000000000000000001000000000000"),
("000000000000100000000000000000000111111111111111111110000000000000000000000000000000000000000011111111111111111111000000000000000000001000000000000"),
("000000000000100000000000000000001111111111111111111111000000000000000000000000000000000000000111111111111111111111100000000000000000001000000000000"),
("000000000000100000000000000000001111111111111111111111100000000000000000000000000000000000001111111111111111111111100000000000000000001000000000000"),
("000000000000100000000000000000011111111111111111111111100000000000000000000000000000000000001111111111111111111111110000000000000000001000000000000"),
("000000000000100000000000000000011111111111111111111111100000000000000000000000000000000000001111111111111111111111110000000000000000001000000000000"),
("000000000000100000000000000000011111111111111111111111100000000000000000000000000000000000011111111111111111111111110000000000000000001000000000000"),
("000000000000100000000000000000011111111111111111111111110000000000000000000000000000000000011111111111111111111111110000000000000000001000000000000"),
("000000000000100000000000000000011111111111111111111111110000000000000000000000000000000000011111111111111111111111110000000000000000001000000000000"),
("000000000000100000000000000000011111111111111111111111110000000000000000000000000000000000011111111111111111111111110000000000000000001000000000000"),
("000000000000100000000000000000011111111111111111111111110000000000000000000000000000000000011111111111111111111111110000000000000000001000000000000"),
("000000000000100000000000000000011111111111111111111111100000000000000000000000000000000000011111111111111111111111110000000000000000001000000000000"),
("000000000000100000000000000000011111111111111111111111100000000000000000000000000000000000001111111111111111111111110000000000000000001000000000000"),
("000000000000100000000000000000011111111111111111111111100000000000000000000000000000000000001111111111111111111111110000000000000000001000000000000"),
("000000000000100000000000000000001111111111111111111111100000000000000000000000000000000000001111111111111111111111100000000000000000001000000000000"),
("000000000000100000000000000000001111111111111111111111000000000000000000000000000000000000000111111111111111111111100000000000000000001000000000000"),
("000000000000100000000000000000000111111111111111111111000000000000000000000000000000000000000111111111111111111111000000000000000000001000000000000"),
("000000000000100000000000000000000111111111111111111110000000000000000000000000000000000000000011111111111111111110000000000000000000001000000000000"),
("000000000000100000000000000000000011111111111111111100000000000000000000000000000000000000000001111111111111111110000000000000000000001000000000000"),
("000000000000100000000000000000000001111111111111111000000000000000000000000000000000000000000000111111111111111000000000000000000000001000000000000"),
("000000000000100000000000000000000000011111111111100000000000000000000000000000000000000000000000001111111111110000000000000000000000001000000000000"),
("000000000000100000000000000000000000000111111110000000000000000000000000000000000000000000000000000011111111000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000111111111000000000000000000000000000000000000000000000000000111111111000000000000000000000000001000000000000"),
("000000000000100000000000000000000000011111111111100000000000000000000000000000000000000000000000011111111111110000000000000000000000001000000000000"),
("000000000000100000000000000000000001111111111111111000000000000000000000000000000000000000000000111111111111111100000000000000000000001000000000000"),
("000000000000100000000000000000000011111111111111111100000000000000000000000000000000000000000001111111111111111110000000000000000000001000000000000"),
("000000000000100000000000000000000111111111111111111110000000000000000000000000000000000000000011111111111111111111000000000000000000001000000000000"),
("000000000000100000000000000000000111111111111111111111000000000000000000000000000000000000000111111111111111111111000000000000000000001000000000000"),
("000000000000100000000000000000001111111111111111111111000000000000000000000000000000000000000111111111111111111111100000000000000000001000000000000"),
("000000000000100000000000000000001111111111111111111111100000000000000000000000000000000000001111111111111111111111100000000000000000001000000000000"),
("000000000000100000000000000000011111111111111111111111100000000000000000000000000000000000001111111111111111111111110000000000000000001000000000000"),
("000000000000100000000000000000011111111111111111111111100000000000000000000000000000000000001111111111111111111111110000000000000000001000000000000"),
("000000000000100000000000000000011111111111111111111111110000000000000000000000000000000000011111111111111111111111110000000000000000001000000000000"),
("000000000000100000000000000000011111111111111111111111110000000000000000000000000000000000011111111111111111111111110000000000000000001000000000000"),
("000000000000100000000000000000011111111111111111111111110000000000000000000000000000000000011111111111111111111111110000000000000000001000000000000"),
("000000000000100000000000000000011111111111111111111111110000000000000000000000000000000000011111111111111111111111110000000000000000001000000000000"),
("000000000000100000000000000000011111111111111111111111110000000000000000000000000000000000011111111111111111111111110000000000000000001000000000000"),
("000000000000100000000000000000011111111111111111111111100000000000000000000000000000000000011111111111111111111111110000000000000000001000000000000"),
("000000000000100000000000000000011111111111111111111111100000000000000000000000000000000000001111111111111111111111110000000000000000001000000000000"),
("000000000000100000000000000000011111111111111111111111100000000000000000000000000000000000001111111111111111111111110000000000000000001000000000000"),
("000000000000100000000000000000001111111111111111111111000000000000000000000000000000000000001111111111111111111111100000000000000000001000000000000"),
("000000000000100000000000000000001111111111111111111111000000000000000000000000000000000000000111111111111111111111100000000000000000001000000000000"),
("000000000000100000000000000000000111111111111111111110000000000000000000000000000000000000000011111111111111111111000000000000000000001000000000000"),
("000000000000100000000000000000000011111111111111111110000000000000000000000000000000000000000011111111111111111110000000000000000000001000000000000"),
("000000000000100000000000000000000001111111111111111100000000000000000000000000000000000000000001111111111111111100000000000000000000001000000000000"),
("000000000000100000000000000000000000111111111111110000000000000000000000000000000000000000000000111111111111111000000000000000000000001000000000000"),
("000000000000100000000000000000000000011111111111100000000000000000000000000000000000000000000000001111111111110000000000000000000000001000000000000"),
("000000000000100000000000000000000000000011111110000000000000000000000000000000000000000000000000000011111110000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000001111000000000000000000000000000000000000000000000000000000000111100000000000000000000000000001000000000000"),
("000000000000100000000000000000000000001111111111000000000000000000000000000000000000000000000000000111111111100000000000000000000000001000000000000"),
("000000000000100000000000000000000000111111111111110000000000000000000000000000000000000000000000011111111111111000000000000000000000001000000000000"),
("000000000000100000000000000000000001111111111111111000000000000000000000000000000000000000000000111111111111111100000000000000000000001000000000000"),
("000000000000100000000000000000000011111111111111111100000000000000000000000000000000000000000001111111111111111110000000000000000000001000000000000"),
("000000000000100000000000000000000111111111111111111110000000000000000000000000000000000000000011111111111111111111000000000000000000001000000000000"),
("000000000000100000000000000000000111111111111111111111000000000000000000000000000000000000000111111111111111111111000000000000000000001000000000000"),
("000000000000100000000000000000001111111111111111111111000000000000000000000000000000000000000111111111111111111111100000000000000000001000000000000"),
("000000000000100000000000000000001111111111111111111111100000000000000000000000000000000000001111111111111111111111100000000000000000001000000000000"),
("000000000000100000000000000000011111111111111111111111100000000000000000000000000000000000001111111111111111111111110000000000000000001000000000000"),
("000000000000100000000000000000011111111111111111111111100000000000000000000000000000000000001111111111111111111111110000000000000000001000000000000"),
("000000000000100000000000000000011111111111111111111111110000000000000000000000000000000000011111111111111111111111110000000000000000001000000000000"),
("000000000000100000000000000000011111111111111111111111110000000000000000000000000000000000011111111111111111111111110000000000000000001000000000000"),
("000000000000100000000000000000011111111111111111111111110000000000000000000000000000000000011111111111111111111111110000000000000000001000000000000"),
("000000000000100000000000000000011111111111111111111111110000000000000000000000000000000000011111111111111111111111110000000000000000001000000000000"),
("000000000000100000000000000000011111111111111111111111110000000000000000000000000000000000011111111111111111111111110000000000000000001000000000000"),
("000000000000100000000000000000011111111111111111111111100000000000000000000000000000000000001111111111111111111111110000000000000000001000000000000"),
("000000000000100000000000000000011111111111111111111111100000000000000000000000000000000000001111111111111111111111110000000000000000001000000000000"),
("000000000000100000000000000000011111111111111111111111100000000000000000000000000000000000001111111111111111111111100000000000000000001000000000000"),
("000000000000100000000000000000001111111111111111111111000000000000000000000000000000000000000111111111111111111111100000000000000000001000000000000"),
("000000000000100000000000000000001111111111111111111111000000000000000000000000000000000000000111111111111111111111000000000000000000001000000000000"),
("000000000000100000000000000000000111111111111111111110000000000000000000000000000000000000000011111111111111111111000000000000000000001000000000000"),
("000000000000100000000000000000000011111111111111111100000000000000000000000000000000000000000001111111111111111110000000000000000000001000000000000"),
("000000000000100000000000000000000001111111111111111000000000000000000000000000000000000000000000111111111111111100000000000000000000001000000000000"),
("000000000000100000000000000000000000111111111111110000000000000000000000000000000000000000000000011111111111111000000000000000000000001000000000000"),
("000000000000100000000000000000000000001111111111000000000000000000000000000000000000000000000000000111111111100000000000000000000000001000000000000"),
("000000000000100000000000000000000000000001111000000000000000000000000000000000000000000000000000000000111100000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000"),
("000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000"),
("000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000")

    );
  
 --define array to hold medium dice bitmaps
 type t_medium_dice_bitmap is array (0 to 49) of std_logic_vector(0 to 48);
	
    --initial display as ZERO
    constant medium_dice_bitmap_0 : t_medium_dice_bitmap := 
    (
("0000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000"),
("0001111111111111111111111111111111111111111111000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001111111111111111111111111111111111111111111000"),
("0000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000")
);
    
    --dice number 1
    constant medium_dice_bitmap_1 : t_medium_dice_bitmap := 
    (
("0000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000"),
("0001111111111111111111111111111111111111111111000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000011000000000000000000001000"),
("0001000000000000000001111110000000000000000001000"),
("0001000000000000000011111111000000000000000001000"),
("0001000000000000000111111111100000000000000001000"),
("0001000000000000000111111111100000000000000001000"),
("0001000000000000000111111111100000000000000001000"),
("0001000000000000000111111111100000000000000001000"),
("0001000000000000000011111111000000000000000001000"),
("0001000000000000000001111110000000000000000001000"),
("0001000000000000000000011000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001111111111111111111111111111111111111111111000"),
("0000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000")
);


--dice number 2
    constant medium_dice_bitmap_2 : t_medium_dice_bitmap := 
    (
("0000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000"),
("0001111111111111111111111111111111111111111111000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000111000000000000000000000000000001000"),
("0001000000001111100000000000000000000000000001000"),
("0001000000011111110000000000000000000000000001000"),
("0001000000111111111000000000000000000000000001000"),
("0001000000111111111000000000000000000000000001000"),
("0001000000111111111000000000000000000000000001000"),
("0001000000111111111000000000000000000000000001000"),
("0001000000011111110000000000000000000000000001000"),
("0001000000001111100000000000000000000000000001000"),
("0001000000000111000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000011100000000001000"),
("0001000000000000000000000000000111110000000001000"),
("0001000000000000000000000000001111111000000001000"),
("0001000000000000000000000000011111111100000001000"),
("0001000000000000000000000000011111111100000001000"),
("0001000000000000000000000000011111111100000001000"),
("0001000000000000000000000000011111111100000001000"),
("0001000000000000000000000000001111111000000001000"),
("0001000000000000000000000000000111110000000001000"),
("0001000000000000000000000000000011100000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001111111111111111111111111111111111111111111000"),
("0000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000")

);


--dice number 3
    constant medium_dice_bitmap_3 : t_medium_dice_bitmap := 
    (
("0000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000"),
("0001111111111111111111111111111111111111111111000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000111000000000000000000000000000001000"),
("0001000000011111110000000000000000000000000001000"),
("0001000000111111110000000000000000000000000001000"),
("0001000000111111111000000000000000000000000001000"),
("0001000001111111111000000000000000000000000001000"),
("0001000001111111111000000000000000000000000001000"),
("0001000000111111111000000000000000000000000001000"),
("0001000000111111110000000000000000000000000001000"),
("0001000000011111100000000000000000000000000001000"),
("0001000000000111000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000001110000000000000000001000"),
("0001000000000000000000111111100000000000000001000"),
("0001000000000000000001111111100000000000000001000"),
("0001000000000000000011111111111000000000000001000"),
("0001000000000000000011111111111000000000000001000"),
("0001000000000000000011111111111000000000000001000"),
("0001000000000000000001111111110000000000000001000"),
("0001000000000000000000111111000000000000000001000"),
("0001000000000000000000011110000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000001111110000001000"),
("0001000000000000000000000000000011111111000001000"),
("0001000000000000000000000000000011111111000001000"),
("0001000000000000000000000000000111111111100001000"),
("0001000000000000000000000000000111111111100001000"),
("0001000000000000000000000000000111111111100001000"),
("0001000000000000000000000000000011111111000001000"),
("0001000000000000000000000000000011111111000001000"),
("0001000000000000000000000000000001111100000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001111111111111111111111111111111111111111111000"),
("0000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000")

);


--dice number 4
    constant medium_dice_bitmap_4 : t_medium_dice_bitmap := 
    (
("0000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000"),
("0001111111111111111111111111111111111111111111000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000111000000000000000001110000000001000"),
("0001000000001111100000000000000011111000000001000"),
("0001000000011111110000000000000111111100000001000"),
("0001000000111111111000000000001111111110000001000"),
("0001000000111111111000000000001111111110000001000"),
("0001000000111111111000000000001111111110000001000"),
("0001000000111111111000000000001111111110000001000"),
("0001000000011111110000000000000111111100000001000"),
("0001000000001111100000000000000011111000000001000"),
("0001000000000111000000000000000001110000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000111000000000000000001110000000001000"),
("0001000000001111100000000000000011111000000001000"),
("0001000000011111110000000000000111111100000001000"),
("0001000000111111111000000000001111111110000001000"),
("0001000000111111111000000000001111111110000001000"),
("0001000000111111111000000000001111111110000001000"),
("0001000000111111111000000000001111111110000001000"),
("0001000000011111110000000000000111111100000001000"),
("0001000000001111100000000000000011111000000001000"),
("0001000000000111000000000000000001110000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001111111111111111111111111111111111111111111000"),
("0000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000")

);


--dice number 5
    constant medium_dice_bitmap_5 : t_medium_dice_bitmap := 
    (
("0000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000"),
("0001111111111111111111111111111111111111111111000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000111000000000000000001110000000001000"),
("0001000000011111110000000000000111111100000001000"),
("0001000000111111110000000000001111111100000001000"),
("0001000000111111111000000000001111111110000001000"),
("0001000000111111111000000000001111111110000001000"),
("0001000000111111111000000000001111111110000001000"),
("0001000000111111110000000000001111111110000001000"),
("0001000000011111110000000000000111111100000001000"),
("0001000000000111000000000000000001110000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000011100000000000000000001000"),
("0001000000000000000000111110000000000000000001000"),
("0001000000000000000001111111000000000000000001000"),
("0001000000000000000011111111100000000000000001000"),
("0001000000000000000011111111100000000000000001000"),
("0001000000000000000011111111100000000000000001000"),
("0001000000000000000011111111100000000000000001000"),
("0001000000000000000001111111000000000000000001000"),
("0001000000000000000000111110000000000000000001000"),
("0001000000000000000000011100000000000000000001000"),
("0001000000000111000000000000000001110000000001000"),
("0001000000001111100000000000000011111000000001000"),
("0001000000011111110000000000000111111100000001000"),
("0001000000111111111000000000001111111110000001000"),
("0001000000111111111000000000001111111110000001000"),
("0001000000111111111000000000001111111110000001000"),
("0001000000111111111000000000001111111110000001000"),
("0001000000011111110000000000000111111100000001000"),
("0001000000001111100000000000000011111000000001000"),
("0001000000000111000000000000000001110000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001111111111111111111111111111111111111111111000"),
("0000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000")

);


--dice number 6
    constant medium_dice_bitmap_6 : t_medium_dice_bitmap := 
    (
("0000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000"),
("0001111111111111111111111111111111111111111111000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000111000000000000000001110000000001000"),
("0001000000001111100000000000000011111000000001000"),
("0001000000011111110000000000000111111100000001000"),
("0001000000111111111000000000001111111110000001000"),
("0001000000111111111000000000001111111110000001000"),
("0001000000111111111000000000001111111110000001000"),
("0001000000111111111000000000001111111110000001000"),
("0001000000011111110000000000000111111100000001000"),
("0001000000001111100000000000000011111000000001000"),
("0001000000000111000000000000000001110000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000111000000000000000001110000000001000"),
("0001000000001111100000000000000011111000000001000"),
("0001000000011111110000000000000111111100000001000"),
("0001000000111111111000000000001111111110000001000"),
("0001000000111111111000000000001111111110000001000"),
("0001000000111111111000000000001111111110000001000"),
("0001000000111111111000000000001111111110000001000"),
("0001000000011111110000000000000111111100000001000"),
("0001000000001111100000000000000011111000000001000"),
("0001000000000111000000000000000001110000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000111000000000000000001110000000001000"),
("0001000000001111100000000000000011111000000001000"),
("0001000000011111110000000000000111111100000001000"),
("0001000000111111111000000000001111111110000001000"),
("0001000000111111111000000000001111111110000001000"),
("0001000000111111111000000000001111111110000001000"),
("0001000000111111111000000000001111111110000001000"),
("0001000000011111110000000000000111111100000001000"),
("0001000000001111100000000000000011111000000001000"),
("0001000000000111000000000000000001110000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001000000000000000000000000000000000000000001000"),
("0001111111111111111111111111111111111111111111000"),
("0000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000")

);


type t_small_dice_bitmap is array (0 to 29) of std_logic_vector(0 to 28);
	
    --dice number 1
    constant small_dice_bitmap_1 : t_small_dice_bitmap := 
    (
("00000000000000000000000000000"),
("00000000000000000000000000000"),
("00111111111111111111111111110"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100000000001110000000000010"),
("00100000000011111000000000010"),
("00100000000011111000000000010"),
("00100000000011111000000000010"),
("00100000000001110000000000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00111111111111111111111111110"),
("00000000000000000000000000000")

);


--dice number 2
    constant small_dice_bitmap_2 : t_small_dice_bitmap := 
    (
("00000000000000000000000000000"),
("00000000000000000000000000000"),
("00111111111111111111111111110"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100001110000000000000000010"),
("00100011111000000000000000010"),
("00100011111000000000000000010"),
("00100011111000000000000000010"),
("00100001110000000000000000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100000000000000001110000010"),
("00100000000000000011111000010"),
("00100000000000000011111000010"),
("00100000000000000011111000010"),
("00100000000000000001110000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00111111111111111111111111110"),
("00000000000000000000000000000")


);


--dice number 3
    constant small_dice_bitmap_3 : t_small_dice_bitmap := 
    (
("00000000000000000000000000000"),
("00000000000000000000000000000"),
("00111111111111111111111111110"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100001110000000000000000010"),
("00100011111000000000000000010"),
("00100011111000000000000000010"),
("00100011111000000000000000010"),
("00100001110000000000000000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100000000001110000000000010"),
("00100000000011111000000000010"),
("00100000000011111000000000010"),
("00100000000011111000000000010"),
("00100000000001110000000000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100000000000000001110000010"),
("00100000000000000011111000010"),
("00100000000000000011111000010"),
("00100000000000000011111000010"),
("00100000000000000001110000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00111111111111111111111111110"),
("00000000000000000000000000000")

);


--dice number 4
    constant small_dice_bitmap_4 : t_small_dice_bitmap := 
    (
("00000000000000000000000000000"),
("00000000000000000000000000000"),
("00111111111111111111111111110"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100001110000000001110000010"),
("00100011111000000011111000010"),
("00100011111000000011111000010"),
("00100011111000000011111000010"),
("00100001110000000001110000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100001110000000001110000010"),
("00100011111000000011111000010"),
("00100011111000000011111000010"),
("00100011111000000011111000010"),
("00100001110000000001110000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00111111111111111111111111110"),
("00000000000000000000000000000")

);


--dice number 5
    constant small_dice_bitmap_5 : t_small_dice_bitmap := 
    (
("00000000000000000000000000000"),
("00000000000000000000000000000"),
("00111111111111111111111111110"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100001110000000001110000010"),
("00100011111000000011111000010"),
("00100011111000000011111000010"),
("00100011111000000011111000010"),
("00100001110000000001110000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100000000001110000000000010"),
("00100000000011111000000000010"),
("00100000000011111000000000010"),
("00100000000011111000000000010"),
("00100000000001110000000000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100001110000000001110000010"),
("00100011111000000011111000010"),
("00100011111000000011111000010"),
("00100011111000000011111000010"),
("00100001110000000001110000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00111111111111111111111111110"),
("00000000000000000000000000000")

);


--dice number 6
    constant small_dice_bitmap_6 : t_small_dice_bitmap := 
    (
("00000000000000000000000000000"),
("00000000000000000000000000000"),
("00111111111111111111111111110"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100001110000000001110000010"),
("00100011111000000011111000010"),
("00100011111000000011111000010"),
("00100011111000000011111000010"),
("00100001110000000001110000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100001110000000001110000010"),
("00100011111000000011111000010"),
("00100011111000000011111000010"),
("00100011111000000011111000010"),
("00100001110000000001110000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100001110000000001110000010"),
("00100011111000000011111000010"),
("00100011111000000011111000010"),
("00100011111000000011111000010"),
("00100001110000000001110000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00100000000000000000000000010"),
("00111111111111111111111111110"),
("00000000000000000000000000000")

);

--CRAPS TABLE 
type t_craps_table_bitmap is array (0 to 432) of std_logic_vector(0 to 639);

constant craps_table_bitmap : t_craps_table_bitmap := 
    (

        ("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000"),
("0000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000"),
("0000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000"),
("0000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000"),
("0000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000"),
("0000000000000000000000000000011111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000000000000000000000000000111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000000000000000000000000000111111110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000000000000000000000000001111111110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000000000000000000000000001111111110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000000000000000000000000011111111110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000000000000000000000000011111011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000000000000000000000000111111011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000000000000000000000000111111011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000000000000000000000001111110011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000000000000000000000001111100011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000000000000000000000011111000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000000000000000000000011111000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000000000000000000000011111000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000000000000000000000111110000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000000000000000000000111110000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000000000000000000001111110000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000000000000000000011111000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000000000000000000011111000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000000000000000000011111000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000000000000000000011110000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000000000000000000111110000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000000000000000001111100000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000000000000000001111100000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000000000000000011111000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000000000000000011111000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000000000000000011111000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000000000000000111111000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000000000000000111110000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000000000000001111100000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000000000000001111100000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000000000000011111000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000000000000011111000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000000000000011111000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000000000000011111000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000000000001111110000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000000000001111100000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000000000001111000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000000000011111000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000000000111111000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000000001111100000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000000001111100000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000000001111100000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000000011111100000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000000011111000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000000111111000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000000111110000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000011000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000111100000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000001111100000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000011111100000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000111111110000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000001111111111000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000011110000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000111000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000111110000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000001111000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000001111100001100000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000111111100000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000011111000000000000000000000000111100000000000000000000000000000000000111111111111110000000000000000000000000000111110000000000000000000000000000000000000000000000000000111111000001100000000000001111100000000000000000000000011110000000000000000000000111111111100000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000001111111100000000000000000000000111110000000000000000000000000000000011111111111111111111111111111100000000000000011111000000000000000000000000000000000000000000000000111111000000000000000000000000111100000000000000000000000000000001111111111111111111110000000000000000000000000111110000000000000000000000000000000000000000000000000000111110000001100000000000001111100000000000000000000000111110000000000000000000011111111111111000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000011111111100000000000000000000000111110000000000000000000000000000000111111111111111111111111111111110000000000000011111000000000000000000000000000000000000000000000001111110000000000000000000000000111100000000000000000000000000000011111111111111111111110000000000000000000000000111110000000000000000000000000000000000000000000000000000111110000001111000000000001111100000000000000000000001111110000000000000000000111111111111111100000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000011111111110000000000000000000000111110000000000000000000000000000000111111111111111111111111111111000000000000000011111000000000000000000000000000000000000000000000001111110000000000000000000000000111100000000000000000000000000001111111111111111111111111110000000000000000000000111110000000000000000000000000000000000000000000000000001111111000001111000000000001111100000000000000001001111111110000000000000000111111111111111111111100000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000111111111110000000000000000000000111110000000000000000000000000000000111111111111111111111111111111000000000000000011111000000000000000000000000000000000000000000000001111110000000000000000000000000111100000000000000000000000000011111111111111111111111111111000000000000000000000111110000000000000000000000000000000000000000000000000001111111100001111000000000001111100000000000000001111111111111000000000000000111111111111111111111110000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000001111111111100000000000000000000000111110000000000000000000000000000001111111111111111111111111111111000000000000000011111000000000000000000000000000000000000000000000000001110000000000000000000000000111100000000000000000000000001111111111111100000111111111111100000000000000000000111110000000000000000000000000000000000000000000000000111111111110001111100000000001111100000000000001111111111111111000000000000011111111111000111111111111000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000011111111111100000000000000000000000111110000000000000000000000000000001111111111111111111111111111111000000000000000011111000000000000000000000000000000000000000000000000001110000000000000000000000000111100000000000000000000000011111111111111000000001111111111110000000000000000000111110000000000000000000000000000000000000000000000000111111111111001111100000011001111100000000000111111111111111110000000000000111111111110000001111111111100000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000011111111111100000000000000000000000111110000000000000000000000000000001111111111111111111111111111111000000000000000011111000000000000000000000000000000000000000000000000001110000000000000000000000000111100000000000000000000000011111111111111000000000111111111111000000000000000000111110000000000000000000000000000000000000000000000000110011111111001111100000011001111100000000000111111111111111110000000000000111111111110000001111111111110000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000011111111111100000000000000000000000111110000000000000000000000000000001111111111111111111111111111111000000000000000011111000000000000000000000000000000000000000000110000001110000000000000000000000000111100000000000000000000000111111111111110000000000111111111111000000000000000000111110000000000000000000000000000000000000000000000111000001111111111111110000011001111100000000111111111111111111111000000000011111111111000000000111111111110000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000001111111111111100000000000000000000000111110000000000000000000000000000111111111111111111111111111111110000000000000000011111000000000000000000000000000000000000000001110000001110000000000000000000000000111100000000000000000000000111111111111100000000000111111111111100000000000000000111110000000000000000000000000000000000000000000000111000000111111111111111000011111111100000111111111111111111111111000000000011111111111100000000111111111111000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000001111111111111100000000000000000000000111110000000000000000000000000000111111111111111111111111111111100000000000000000011111000000000000000000000000000000000000000001110000001110000000000000000000000000111100000000000000000000001111111111111000000000000011111111111100000000000000000111110000000000000000000000000000000000000000000001111100000111111111000011000011111111100001111111111111111111111110000000000011111111111100000000111111111111000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000011111111111111100000000000000000000000111110000000000000000000000000000111111111111111111111111111111100000000000000000011111000000000000000000000000000000000000000111110000001100000000000000000000000000111100000000000000000000011111111111111000000000000001111111111110000000000000000111110000000000000000000000000000000000000000000111110000000111111111000000000011111111100111111111111111111111111111000000001111111111111000000000001111111111100000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000111111111111111100000000000000000000000111110000000000000000000000000000111111111111111111111111111111100000000000000000011111000000000000000000000000000000000000001111111110001100000000000000000000000000111100000000000000000000011111111111111000000000000001111111111111000000000000000111110000000000000000000000000000000000000000001111110000000011111111100000000011111111100111111111111111111111111111000000001111111111111000000000001111111111100000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000111111111111111100000000000000000000000111110000000000000000000000000001111111111111111111111111111111110000000000000000011111000000000000000000000000000000000000001111111110001110000000000000000000000000111100000000000000000000011111111111111000000000000001111111111111000000000000000111110000000000000000000000000000000000000000001111110000000001111111100000000011111111100111000000011111111111111111000000001111111111110000000000001111111111110000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000001111111111111111100000000000000000000000111110000000000000000000000000011111111111111111111111011111110000000000000000000011111000000000000000000000000000000000000011111111111111110000000000000000000000000111100000000000000000000011111111111111000000000000001111111111111000000000000000111110000000000000000000000000000000000000000011111110000000001111111100000001111111111100000000000001111111111111110000000011111111111110000000000001111111111100000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000011111111111111111100000000000000000000000111110000000000000000000000000011111100000000000000000000000000000000000000000000011111000000000000000000000000000000000000111111111111111111000000000000000000000000111100000000000000000000011111111111111000000000000001111111111111000000000000000111110000000000000000000000000000000000000000011111111000000000111111110000001111111111100000000000001111111111111110000000011111111111110000000000001111111111111000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000111111111111111111110000000000000000000000111110000000000000000000000000011111100000000000000000000000000000000000000000000011111000000000000000000000000000000000001111111111111111111100000000000000000000000111100000000000000000000011111111111111100000000000001111111111111000000000000000111110000000000000000000000000000000000000000000000111100000000011111111000001111001111100000000000001111111111111111000000011111111111110000000000001111111111111000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000001111111111111111111100000000000000000000000111110000000000000000000000000111110000000000000000000000000000000000000000000000011111000000000000000000000000000000000111110001111111111111111110000000000000000000111100000000000000000000011111111111111110000000000001111111111111000000000000000111110000000000000000000000000000000000000000000000111100000000011111111000001110001111100000000000001111111111111110000000011111111111110000000000001111111111111000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000001111111111111111111100000000000000000000000111110000000000000000000000000111110000000000000000000000000000000000000000000000011111000000000000000000000000000000001111110000011111111111111111010000000000000000111100000000000000000000011111111111111110000000000001111111111111000000000000000111110000000000000000000000000000000000000000000000011110000000011111111100011100001111100000000000001111111111111110000000111111111111110000000000001111111111111100011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000001111111111111111111100000000000000000000000111110000000000000000000000000111110000000000000000000000000000000000000000000000011111000000000000000000000000000000001110000000001111111111111111111011000000000000111100000000000000000000011111111111111111000000000001111111111111000000000000000111110000000000000000000000000000000000000000000000001110000000001111111110011000001111100000000000001111111111111111000000111111111111110000000000001111111111111100011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000111111011111111111111100000000000000000000000111110000000000000000000000001111111111110000000000000000000000000000000000000000011111000000000000000000000000000000011110000000000000011111111111111111110000000000111100000000000000000000011111111111111111100000000001111111111110000000000000000111110000000000000000000000000000000000000000000000000110000000000111111111111000001111100000000000001111111111111110000000111111111111110000000000001111111111111100011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000111110011111111111111100000000000000000000000111110000000000000000000000001111111111111101100000000000000000000000000000000000011111000000000000000000000000000000111110000000000000001111111111111111110000000000111100000000000000000000011111111111111111110000000011111111111100000000000000000111110000000000000000000000000000000000000100000000000110000000000011111111111000001111100000000000001111111111111110000001111111111111110000000000001111111111111100011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000001111110011111111111111100000000000000000000000111110000000000000000000000001111111111111111111111000000000000000000000000000000011111000000000000000000000000000001111111000000000000001110011111111111000000000000111100000000000000000000001111111111111111110000000011111111111100000000000000000111110000000000000000000000000000000000111110000000000011100000000001111111100000001111100000000000001111111111111111000001111111111111110000000000001111111111111110011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000001111100011111111111111100000000000000000000000111110000000000000000000000011111111111111111111111110000000000000000000000000000011111000000000000000000000000000011111111100000000000001110001111111111000000000000111100000000000000000000011111111111111111111100000111111111111100000000000000000111110000000000000000000000000000000011111111111000000001110000000001111111100000001111100000000000001111111111111111000001111111111111110000000000001111111111111100011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000011111000111111111111111100000000000000000000000111110000000000000000000000011111111111111111111111110000000000000000000000000000011111000000000000000000000000000111111111100000000000001110000011111111000000000000111100000000000000000000011111111111111111111110000111111111111000000000000000000111110000000000000000000000000000000011111111111001000001110000000001111111000000001111100000000000001111111111111110000001111111111111110000000000011111111111111100011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000111110000011111111111111100000000000000000000000111110000000000000000000000111111111111111111111111111111000000000000000000000000011111000000000000000000000000000110111111110000000000001111000001111100000000000000111100000000000000000000001111111111111111111111100111111111100000000000000000000111110000000000000000000000000000000111111111111111111111111000000000111110000000001111100000000000001111111111111111000001111111111111110000000000001111111111111110011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000111110000011111111111111100000000000000000000000111110000000000000000000000111111111111111111111111111111100000000000000000000000011111000000000000000000000000000110111111110000000000001110000000111000000000000000111100000000000000000000001111111111111111111111111111111111100000000000000000000111110000000000000000000000000000011111111111111111111111111100000001111100000000001111100000000000001111111111111111000011111111111111110000000000001111111111111111011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000001111100000011111111111111100000000000000000000000111110000000000000000000000111111111111111111111111111111100000000000000000000000011111000000000000000000000000000100011111110000000000001100000000111000000000000000111100000000000000000000001111111111111111111111111111111110000000000000000000000111110000000000000000000000000000011111111111111111111111111100000001111000000000001111100000000000001111111111111110000011111111111111110000000000001111111111111111011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000111111000000011111111111111110000000000000000000000111110000000000000000000000111111111111111111111111111111111000000000000000000000011111000000000000000000000000000000001111111100000000001111000000000000000000000000111100000000000000000000000011111111111111111111111111111100000000000000000000000111110000000000000000000000000000000000111111111111111111111110000000100000000000001111100000000000001111111111111111000011111111111111110000000000001111111111111111011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000111110000000011111111111111110000000000000000000000111110000000000000000000011111111111111111111111111111111111110000000000000000000011111000000000000000000000110000000001111111100000000001110000000000000000000000000111100000000000000000000000011111111111111111111111111111100000000000000000000000111110000000000000000000000000001100000111111111111111111111110000000000000000000001111100000000000001111111111111111000011111111111111110000000000001111111111111111011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000111110000000111111111111111100000000000000000000000111110000000000000000000011111111111111111111111111111111111111000000000000000000011111000000000000000000000111000000000111111100000000001110000000000000000000000000111100000000000000000000000000111111111111111111111111100000000000000000000000000111110000000000000000000000000011100000011110000111111111111110000000000000000000001111100000000000001111111111111110000011111111111111110000000000001111111111111111011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000001111100000000011111111111111100000000000000000000000111110000000000000000000011111111111111111111111111111111111111000000000000000000011111000000000000000000011111100000000011111110000000001110000000000000000000000000111100000000000000000000000000011111111111111111111111110000000000000000000000000111110000000000000000000000000011100000000110000011111111111111100000000000000000001111100000000000001111111111111111000011111111111111110000000000001111111111111111011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000011111100000000011111111111111100000000000000000000000111110000000000000000000011111111111111111111111111111111111111000000000000000000011111000000000000000000111111110000000011111110000000001111100000000000000000000000111100000000000000000000000000011111111111111111111111111000000000000000000000000111110000000000000000000000000011100000000111000001001111111111100000000000000000001111100000000000001111111111111111000011111111111111110000000000001111111111111111011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000111110000000000011111111111111100000000000000000000000111110000000000000000000111111111111111111111111111111111111111100000000000000000011111000000000000000011111111111000000001111110000000001111111000000000000000000000111100000000000000000000000000000011111111111111111111111100000000000000000000000111110000000000000000000000001111000000000111000000000010111111100000000000000000001111100000000000001111111111111110000011111111111111110000000000111111111111111111011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000111110000000000001111111111111110000000000000000000000111110000000000000000000011111111111111111111111111111111111111110000000000000000011111000000000000000011111111111000000000111111100000001111100000000000000000000000111100000000000000000000000000000001111111111111111111111111000000000000000000000111110000000000000000000000011111100000000011000000000000001111000000000000000000001111100000000000001111111111111111000011111111111111110000000000001111111111111111011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000111110000000000001111111111111110000000000000000000000111110000000000000000000000000000000111111111111111111111111111111000000000000000011111000000000000000111111111111000000000111111110000001111100000000000000000000000111100000000000000000000000000000000111111111111111111111111100000000000000000000111110000000000000000000000011111100000000011100000000000000110000000000000000000001111100000000000001111111111111111000011111111111111110000000000001111111111111111011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000011111100000000000111111111111111100000000000000000000000111110000000000000000000000000000000000000111111111111111111111111000000000000000011111000000000000011111000000111100000000111111110000011111000000000000000000000000111100000000000000000000000000000001111111111111111111111111100000000000000000000111110000000000000000000001111111110000000001110000000000000000000000000000000000001111100000000000001111111111111110000011111111111111110000000000001111111111111111011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000111111000000000000011111111111111100000000000000000000000111110000000000000000000000000000000000000011111111111111111111111000000000000000011111000000000000011110000000011100000000111111110000011110000000000000000000000000111100000000000000000000000000000111111111111111111111111111111000000000000000000111110000000000000000000011111111111000000000111000000000000000000000000000000000001111100000000000001111111111111110000011111111111111110000000000001111111111111111011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000111110000000000000011111111111111100000000000000000000000111110000000000000000000000000000000000000001111111111111111111111000000000000000011111000000000000011100000000001100000000011111110000011100000000000000000000000000111100000000000000000000000000000111111111111111111111111111111000000000000000000111110000000000000000000011111111111000000000111000000000000000000000000000000000001111100000000000001111111111111111000011111111111111110000000000001111111111111111011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000111110000000000000111111111111111100000000000000000000000111110000000000000000000000000000000000000000001111111111111111111000000000000000011111000000000000011100000000000000000000000111111101100000000000000000000000000000111100000000000000000000000000011111111100111111111111111111111100000000000000000111110000000000000000000011101111111000000000111000000000000000000000000000000000001111100000000000001111111111111110000011111111111111110000000000011111111111111111011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000011111110000000000000001111111111111110000000000000000000000111110000000000000000000000000000000000000000000011111111111111111110000000000000011111000000000000111100000000000000000000000111111111100000000000000000000000000000111100000000000000000000000011111111111000011111111111111111111100000000000000000111110000000000000000011000001111111110000000011110000000000000000000000000000000001111100000000000001111111111111111000011111111111111110000000000001111111111111111011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000011111000000000000000001111111111111110000000000000000000000111110000000000000000000000000000000000000000000001111111111111111110000000000000011111000000000001111110000000000000000000000111111111100000000000000000000000000000111100000000000000000000000011111111110000001111111111111111111100000000000000000111110000000000000000111100000011111110000000011110000000000000000000000000000000001111100000000000001111111111111111000011111111111111110000000000001111111111111111011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000111111111111111111111111111111111111111111000000000000000000111110000000000000000000000000000000000000000000000001111111111111110000000000000011111000000000000111111111100111111100000000001111110000000000000000000000000000000111100000000000000000000001111111111110000000111111111111111111111000000000000000111110000000000000001111000000011111110000000000111001000000000000000000000000000001111100000000000001111111111111110000011111111111111110000000000001111111111111111011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000111111111111111111111111111111111111111111110000000000000000111110000000000000000000000000000000000000000000000001111111111111110000000000000011111000000000000011111111111111111111110000001111110000000000000000000000000000000111100000000000000000000001111111111110000000011111111111111111111000000000000000111110000000000000011111100000011111111000000000111111100000000000000000000000000001111100000000000001111111111111111000011111111111111110000000000001111111111111111011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000111111111111111111111111111111111111111111110000000000000000111110000000000000000000000000000000000000000000000001111111111111110000000000000011111000000000000011111111111111111111110000001111100000000000000000000000000000000111100000000000000000000001111111111100000000001111111111111111111100000000000000111110000000000000111111100000001111111100000000111111110000000000000000000000000001111100000000000001111111111111111000011111111111111110000000000001111111111111110011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000111111111111111111111111111111111111111111110000000000000000111110000000000000000000000000000000000000000000000000011111111111110000000000000011111000000000000011111111111111111111110000001110000000000000000000000000000000000111100000000000000000000011111111111100000000000111111111111111111100000000000000111110000000000001111111000000001111111110000000011111000000000000000000000000000001111100000000000001111111111111110000001111111111111110000000000001111111111111100011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000111111111111111111111111111111111111111111110000000000000000111110000000000000000000000000000000000000000000000000011111111111110000000000000011111000000000000011111111111111111111111000111110000000000000000000000000000000000111100000000000000000000011111111111000000000000011111111111111111100000000000000111110000000000001111111100000000111111110000000001111000000000000000000000000000001111100000000000001111111111111110000001111111111111110000000000001111111111111100011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000111111111111111111111111111111111111111111110000000000000000111110000000000000000000000000000000000000000000000000001111111111110000000000000011111000000000000001111111111111111111111100111100000000000000000000000000000000000111100000000000000000000011111111111000000000000001111111111111111100000000000000111110000000000001101111100000000011111110000000001110000000000000000000000000000001111100000000000001111111111111111000001111111111111110000000000001111111111111100011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000111111111111111111111111111111111111111111110000000000000000111110000000000000000000000000000000000000000000000000001111111111110000000000000011111000000000000000011111111111111111111100110000000000000000000000000000000000000111100000000000000000001111111111111000000000000001111111111111111100000000000000111110000000000001100111100000000011111111000000011100000000000000000000000000000001111100000000000001111111111111110000001111111111111110000000000011111111111111100011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000111111111111111111111111111111111111111111110000000000000000111110000000000000000000000000000000000000000000000000001111111111110000000000000011111000000000000000011111111111111111111100110000000000000000000000000000000000000111100000000000000000001111111111111000000000000001111111111111111100000000000000111110000000000000000011100000000011111111000000011100000000000000000000000000000001111100000000000001111111111111110000001111111111111110000000000011111111111111100011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000111111111111111111111111111111111111111111110000000000000000111110000000000000000000000000000000000000000000000000000111111111110000000000000011111000000000000000000000000000000011111100000000000000000000000000000000000000000111100000000000000000001111111111111000000000000000111111111111111100000000000000111110000000000000000001111000000000111111100000001100000000000000000000000000000001111100000000000001111111111111111000000111111111111110000000000001111111111111100011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000111111111111111111111111111111111111111111110000000000000000111110000000000000000000000000000000000000000000000000000011111111000000000000000011111000000000000000000000000000000001111100000000000000000000000000000000000000000111100000000000000000001111111111111000000000000000111111111111111100000000000000111110000000000000000001111000000000011111110110000000000000000000000000000000000001111100000000000001111111111111111000000011111111111110000000000001111111111111000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000111111111111111111111111111111111111111111100000000000000000111110000000000000000000000000000000000000000000000000000011111111000000000000000011111000000000000000000000000000000001111100000000000000000000000000000000000000000111100000000000000000001111111111111000000000000000111111111111111100000000000000111110000000000000000001111000000000011111110111000000000000000000000000000000000001111100000000000001111111111111110000000011111111111110000000000011111111111111000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000011111111111111110000000000000000000000111110000000000000000000000000000000000000000000000000000011111111000000000000000011111000000000000000000000000000000000111100000000000000000000000000000000000000000111100000000000000000001111111111111000000000000000111111111111111100000000000000111110000000000000000000011100000000011111111111100000000000000000000000000000000001111100000000000001111111111111111000000011111111111110000000000001111111111111000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000011111111111111100000000000000000000000111110000000000000000000000011011000000000000000000000000011111111000000000000000011111000000000000000000000000000000000111000000000000000000000000000000000000000000111100000000000000000001111111111111000000000000000111111111111111100000000000000111110000111111100000000011110000000011111111110000000000000000000000000000000000001111100000000000001111111111111111000000011111111111110000000000001111111111111000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000011111111111111100000000000000000000000111110000000000000000000000111111000000000000000000000000011111111000000000000000011111000000000000000000011000000000011110000000000000000000000000000000000000000000111100000000000000000001111111111111000000000000000111111111111111100000000000000111110000111111111100000011111000000011111111110000000000000000000000000000000000001111100000000000001111111111111110000000011111111111110000000000001111111111100000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000011111111111111110000000000000000000000111110000000000000000000011111111111000000000000000000000011111110000000000000000011111000000000000000000011111000011111000000000000000000000000000000000000000000000111100000000000000000000111111111111000000000000000011111111111111000000000000000111110011111111111111111001111000000000111111000000000000000000000000000000000000001111100000000000001111111111111111000000001111111111110000000000001111111111110000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000011111111111111110000000000000000000000111110000000000000000000111111111111110000000000000000000011111100000000000000000011111000000000000000000011111111111111000000000000000000000000000000000000000000000111100000000000000000000011111111111000000000000000111111111111111000000000000000111110111111111111111111111111000000000111111000000000000000000000000000000000000001111100000000000001111111111111110000000000111111111111000000000001111111111100000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000111111111111111100000000000000000000000111110000000000000000000111111111111110000000000000000000011111100000000000000000011111000000000000000000000111111111110000000000000000000000000000000000000000000000111100000000000000000000011111111111000000000000000111111111111100000000000000000111110111111111111111111111011000000001111100000000000000000000000000000000000000001111100000000000001111111111111110000000000111111111111000000000001111111111100000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000001111111111111100000000000000000000000111110000000000000000000111111111111111100000000000000000111111000000000000000000011111000000000000000000000111111111000000000000000000000000000000000000000000000000111100000000000000000000011111111111000000000000000111111111111100000000000000000111110010111111111111111111111100000000111000000000000000000000000000000000000000001111100000000000001111111111111111000000000011111111111100000000111111111111000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000011111111111111100000000000000000000000111110000000000000000000111111111111111110000000000000001111111000000000000000000011111000000000000000000000111111110000000000000000000000000000000000000000000000000111100000000000000000000011111111111110000000000001111111111111100000000000000000111110011111111111111111111111100000000111000000000000000000000000000000000000000001111100000000000001111111111111110000000000011111111111100000000111111111111000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000011111111111111100000000000000000000000111110000000000000000000111111111111111111100000000000001111100000000000000000000011111000000000000000000000011111100000000000000000000000000000000000000000000000000111100000000000000000000001111111111110000000000001111111111111000000000000000000111110000111110001111111111111110000011100000000000000000000000000000000000000000001111100000000000001111111111111110000000000011111111111000000000111111111110000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000011111111111111110000000000000000000000111110000000000000000000011111111111111111110000000000011111000000000000000000000011111000000000000000000000001111000000000000000000000000000000000000000000000000000111100000000000000000000000111111111111000000000111111111111110000000000000000000111110000011110000001111111111111100000000000000000000000000000000000000000000000001111100000000000001111111111111111000000000000111111111110000001111111111100000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000011111111111111110000000000000000000000111110000000000000000000011111111111111111111010000001111111000000000000000000000011111000000000000000000000000111000000000000000000000000000000000000000000000000000111100000000000000000000000111111111111110000001111111111111100000000000000000000111110000001110000001111111111111100000000000000000000000000000000000000000000000001111100000000000011111111111111111000000000000111111111111000001111111111100000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000011111111111111100000000000000000000000111110000000000000000000011111111111111111111110000011111100000000000000000000000011111000000000000000000000000100000000000000000000000000000000000000000000000000000111100000000000000000000000001111111111111000001111111111111000000000000000000000111110000000111100000010011111111100000000000000000000000000000000000000000000000001111100000000000111111111111111111100000000000011111111111000111111111110000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000011111111111111100000000000000000000000111110000000000000000000001111111111111111111111111111111100000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000111111111111111111111111111110000000000000000000000111110000000111100000000000011111111000000000000000000000000000000000000000000000001111100000001111111111111111111111111000000000000111111111111111111111100000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000011111111111111100000000000000000000000111110000000000000000000000111111111111111111111111111100000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000011111111111111111111111111100000000000000000000000111110000000011100000000000011111111000000000000000000000000000000000000000000000001111100001111111111111111111111111111111000000000111111111111111111111100000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000011111111111111100000000000000000000000111110000000000000000000000000111111111111111111111110000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000111111111111111111111100000000000000000000000000111110000000001111000000000000001111000000000000000000000000000000000000000000000001111100111111111111111111111111111111111111000000000111111111111111100000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000001111111111111000000000000000000000000111110000000000000000000000000111111111111111111111100000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000011111111111111111111100000000000000000000000000111110000000001111000000000000000000000000000000000000000000000000000000000000000001111100111111111111111111111111111111111111000000000111111111111110000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000111111111111110000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000001111111111110000000000000000000000000000000111110000000000111100000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000111111111100000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000111100000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000111110000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000001110000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000111000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000111000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000111100000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000001111100000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000001111100000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000001111000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000001110000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000001110000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000001110000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000001000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000011111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000"),
("0000001111100000000000000000000011110000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111100000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000001111110000000000000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000111110000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000111111000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000111111000000000000000000000000000001111111111101101100000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000111111000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000011111000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000011111100000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000011111100000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000011111100000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000011111100000000000000000000000000000000000000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000001111111111100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000001111111111111111111011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000001111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000001111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000011111111111111111111111111100000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000")
);
  


  --CRAPS TABLE 
type t_dot is array (0 to 49) of std_logic_vector(0 to 49);

constant dot : t_dot := 
(
("00000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000"),
("00000000000000000000001111110000000000000000000000"),
("00000000000000000000111111111100000000000000000000"),
("00000000000000000011111111111111000000000000000000"),
("00000000000000000111111111111111100000000000000000"),
("00000000000000001111111111111111110000000000000000"),
("00000000000000011111111111111111111000000000000000"),
("00000000000000111111111111111111111100000000000000"),
("00000000000001111111111111111111111110000000000000"),
("00000000000011111111111111111111111111000000000000"),
("00000000000111111111111111111111111111100000000000"),
("00000000001111111111111111111111111111110000000000"),
("00000000011111111111111111111111111111111000000000"),
("00000000111111111111111111111111111111111100000000"),
("00000001111111111111111111111111111111111110000000"),
("00000011111111111111111111111111111111111111000000"),
("00000011111111111111111111111111111111111111000000"),
("00000111111111111111111111111111111111111111100000"),
("00001111111111111111111111111111111111111111110000"),
("00001111111111111111111111111111111111111111110000"),
("00011111111111111111111111111111111111111111111000"),
("00011111111111111111111111111111111111111111111000"),
("00111111111111111111111111111111111111111111111100"),
("00111111111111111111111111111111111111111111111100"),
("00111111111111111111111111111111111111111111111100"),--middle
("00111111111111111111111111111111111111111111111100"),
("00111111111111111111111111111111111111111111111100"),
("00111111111111111111111111111111111111111111111100"),
("00011111111111111111111111111111111111111111111000"),
("00001111111111111111111111111111111111111111110000"),
("00001111111111111111111111111111111111111111100000"),
("00000111111111111111111111111111111111111111100000"),
("00000011111111111111111111111111111111111111000000"),
("00000011111111111111111111111111111111111111000000"),
("00000001111111111111111111111111111111111110000000"),
("00000000111111111111111111111111111111111100000000"),
("00000000011111111111111111111111111111111000000000"),
("00000000001111111111111111111111111111110000000000"),
("00000000000111111111111111111111111111100000000000"),
("00000000000011111111111111111111111111000000000000"),
("00000000000000111111111111111111111100000000000000"),
("00000000000000011111111111111111111000000000000000"),
("00000000000000001111111111111111110000000000000000"),
("00000000000000000111111111111111100000000000000000"),
("00000000000000000011111111111111000000000000000000"),
("00000000000000000000111111111100000000000000000000"),
("00000000000000000000001111110000000000000000000000"),
("00000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000")

);
  

  -----------------------------------------------------------------------------
  -- Numeric bit patterns for output to VGA for scorekeeping
  -----------------------------------------------------------------------------
  


  -----------------------------------------------------------------------------
  -- Component Declarations
  -----------------------------------------------------------------------------
  

  -----------------------------------------------------------------------------
  -- Function Declarations
  -----------------------------------------------------------------------------


    

  
end package bitmaps_pkg;  

package body bitmaps_pkg is


    
end package body bitmaps_pkg;




